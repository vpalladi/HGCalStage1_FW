------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 2.6
--  \   \         Application : 7 Series FPGAs Transceivers Wizard 
--  /   /         Filename : xilinx_gth_16b_5g_cpll_exdes.vhd
-- /___/   /\      
-- \   \  /  \ 
--  \___\/\___\
--
--
-- Module xilinx_gth_16b_5g_cpll_exdes
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

--***********************************Entity Declaration************************

entity xilinx_gth_16b_5g_cpll_exdes is
generic
(
    EXAMPLE_CONFIG_INDEPENDENT_LANES        : integer   := 1;
    STABLE_CLOCK_PERIOD                     : integer   := 32;    --Period of the stable clock driving this state-machine, unit is [ns]
    EXAMPLE_LANE_WITH_START_CHAR            : integer   := 0;    -- specifies lane with unique start frame ch
    EXAMPLE_WORDS_IN_BRAM                   : integer   := 512;  -- specifies amount of data in BRAM
    EXAMPLE_SIM_GTRESET_SPEEDUP             : string    := "TRUE";    -- simulation setting for GT SecureIP model
    EXAMPLE_SIMULATION                      : integer   := 0;             -- Set to 1 for simulation
    EXAMPLE_USE_CHIPSCOPE                   : integer   := 0           -- Set to 1 to use Chipscope to drive resets
);
port
(
    Q7_CLK0_GTREFCLK_PAD_N_IN               : in   std_logic;
    Q7_CLK0_GTREFCLK_PAD_P_IN               : in   std_logic;
    DRP_CLK_IN                              : in   std_logic;
    GTTX_RESET_IN                           : in   std_logic;
    GTRX_RESET_IN                           : in   std_logic;
    CPLL_RESET_IN                           : in   std_logic; 
    QPLL_RESET_IN                           : in   std_logic;
    TRACK_DATA_OUT                          : out  std_logic;
    RXN_IN                                  : in   std_logic_vector(3 downto 0);
    RXP_IN                                  : in   std_logic_vector(3 downto 0);
    TXN_OUT                                 : out  std_logic_vector(3 downto 0);
    TXP_OUT                                 : out  std_logic_vector(3 downto 0)
);


end xilinx_gth_16b_5g_cpll_exdes;
    
architecture RTL of xilinx_gth_16b_5g_cpll_exdes is
    attribute CORE_GENERATION_INFO : string;
    attribute CORE_GENERATION_INFO of RTL : architecture is "xilinx_gth_16b_5g_cpll,gtwizard_v2_6,{protocol_file=Start_from_scratch}";

--**************************Component Declarations*****************************

component xilinx_gth_16b_5g_cpll_init
generic
(
    -- Simulation attributes
    EXAMPLE_SIM_GTRESET_SPEEDUP    : string    := "FALSE";    -- Set to 1 to speed up sim reset
    EXAMPLE_SIMULATION             : integer   := 0;          -- Set to 1 for simulation
    STABLE_CLOCK_PERIOD            : integer   := 32;    --Period of the stable clock driving this state-machine, unit is [ns]
    EXAMPLE_USE_CHIPSCOPE          : integer   := 0           -- Set to 1 to use Chipscope to drive resets
);
port
(
    SYSCLK_IN                               : in   std_logic;
    SOFT_RESET_IN                           : in   std_logic;
    DONT_RESET_ON_DATA_ERROR_IN             : in   std_logic;
    GT0_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_DATA_VALID_IN                       : in   std_logic;
    GT1_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_DATA_VALID_IN                       : in   std_logic;
    GT2_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_DATA_VALID_IN                       : in   std_logic;
    GT3_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT3_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT3_DATA_VALID_IN                       : in   std_logic;

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT0  (X1Y32)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    GT0_CPLLFBCLKLOST_OUT                   : out  std_logic;
    GT0_CPLLLOCK_OUT                        : out  std_logic;
    GT0_CPLLLOCKDETCLK_IN                   : in   std_logic;
    GT0_CPLLRESET_IN                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    GT0_GTREFCLK0_IN                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    GT0_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT0_DRPCLK_IN                           : in   std_logic;
    GT0_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT0_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT0_DRPEN_IN                            : in   std_logic;
    GT0_DRPRDY_OUT                          : out  std_logic;
    GT0_DRPWE_IN                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    GT0_LOOPBACK_IN                         : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    GT0_RXUSERRDY_IN                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    GT0_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    GT0_RXCDRLOCK_OUT                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    GT0_RXUSRCLK_IN                         : in   std_logic;
    GT0_RXUSRCLK2_IN                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    GT0_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    ------------------- Receive Ports - Pattern Checker Ports ------------------
    GT0_RXPRBSERR_OUT                       : out  std_logic;
    GT0_RXPRBSSEL_IN                        : in   std_logic_vector(2 downto 0);
    ------------------- Receive Ports - Pattern Checker ports ------------------
    GT0_RXPRBSCNTRESET_IN                   : in   std_logic;
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    GT0_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT0_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GT0_GTHRXN_IN                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    GT0_RXBYTEISALIGNED_OUT                 : out  std_logic;
    GT0_RXCOMMADET_OUT                      : out  std_logic;
    GT0_RXMCOMMAALIGNEN_IN                  : in   std_logic;
    GT0_RXPCOMMAALIGNEN_IN                  : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    GT0_RXOUTCLK_OUT                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GT0_GTRXRESET_IN                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    GT0_RXPOLARITY_IN                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    GT0_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT0_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    GT0_GTHRXP_IN                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    GT0_RXRESETDONE_OUT                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GT0_GTTXRESET_IN                        : in   std_logic;
    GT0_TXUSERRDY_IN                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    GT0_TXUSRCLK_IN                         : in   std_logic;
    GT0_TXUSRCLK2_IN                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GT0_TXDATA_IN                           : in   std_logic_vector(15 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GT0_GTHTXN_OUT                          : out  std_logic;
    GT0_GTHTXP_OUT                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    GT0_TXOUTCLK_OUT                        : out  std_logic;
    GT0_TXOUTCLKFABRIC_OUT                  : out  std_logic;
    GT0_TXOUTCLKPCS_OUT                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    GT0_TXRESETDONE_OUT                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    GT0_TXPOLARITY_IN                       : in   std_logic;
    ------------------ Transmit Ports - pattern Generator Ports ----------------
    GT0_TXPRBSSEL_IN                        : in   std_logic_vector(2 downto 0);
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    GT0_TXCHARISK_IN                        : in   std_logic_vector(1 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT1  (X1Y33)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    GT1_CPLLFBCLKLOST_OUT                   : out  std_logic;
    GT1_CPLLLOCK_OUT                        : out  std_logic;
    GT1_CPLLLOCKDETCLK_IN                   : in   std_logic;
    GT1_CPLLRESET_IN                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    GT1_GTREFCLK0_IN                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    GT1_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT1_DRPCLK_IN                           : in   std_logic;
    GT1_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT1_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT1_DRPEN_IN                            : in   std_logic;
    GT1_DRPRDY_OUT                          : out  std_logic;
    GT1_DRPWE_IN                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    GT1_LOOPBACK_IN                         : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    GT1_RXUSERRDY_IN                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    GT1_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    GT1_RXCDRLOCK_OUT                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    GT1_RXUSRCLK_IN                         : in   std_logic;
    GT1_RXUSRCLK2_IN                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    GT1_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    ------------------- Receive Ports - Pattern Checker Ports ------------------
    GT1_RXPRBSERR_OUT                       : out  std_logic;
    GT1_RXPRBSSEL_IN                        : in   std_logic_vector(2 downto 0);
    ------------------- Receive Ports - Pattern Checker ports ------------------
    GT1_RXPRBSCNTRESET_IN                   : in   std_logic;
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    GT1_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT1_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GT1_GTHRXN_IN                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    GT1_RXBYTEISALIGNED_OUT                 : out  std_logic;
    GT1_RXCOMMADET_OUT                      : out  std_logic;
    GT1_RXMCOMMAALIGNEN_IN                  : in   std_logic;
    GT1_RXPCOMMAALIGNEN_IN                  : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    GT1_RXOUTCLK_OUT                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GT1_GTRXRESET_IN                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    GT1_RXPOLARITY_IN                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    GT1_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT1_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    GT1_GTHRXP_IN                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    GT1_RXRESETDONE_OUT                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GT1_GTTXRESET_IN                        : in   std_logic;
    GT1_TXUSERRDY_IN                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    GT1_TXUSRCLK_IN                         : in   std_logic;
    GT1_TXUSRCLK2_IN                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GT1_TXDATA_IN                           : in   std_logic_vector(15 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GT1_GTHTXN_OUT                          : out  std_logic;
    GT1_GTHTXP_OUT                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    GT1_TXOUTCLK_OUT                        : out  std_logic;
    GT1_TXOUTCLKFABRIC_OUT                  : out  std_logic;
    GT1_TXOUTCLKPCS_OUT                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    GT1_TXRESETDONE_OUT                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    GT1_TXPOLARITY_IN                       : in   std_logic;
    ------------------ Transmit Ports - pattern Generator Ports ----------------
    GT1_TXPRBSSEL_IN                        : in   std_logic_vector(2 downto 0);
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    GT1_TXCHARISK_IN                        : in   std_logic_vector(1 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT2  (X1Y34)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    GT2_CPLLFBCLKLOST_OUT                   : out  std_logic;
    GT2_CPLLLOCK_OUT                        : out  std_logic;
    GT2_CPLLLOCKDETCLK_IN                   : in   std_logic;
    GT2_CPLLRESET_IN                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    GT2_GTREFCLK0_IN                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    GT2_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT2_DRPCLK_IN                           : in   std_logic;
    GT2_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT2_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT2_DRPEN_IN                            : in   std_logic;
    GT2_DRPRDY_OUT                          : out  std_logic;
    GT2_DRPWE_IN                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    GT2_LOOPBACK_IN                         : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    GT2_RXUSERRDY_IN                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    GT2_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    GT2_RXCDRLOCK_OUT                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    GT2_RXUSRCLK_IN                         : in   std_logic;
    GT2_RXUSRCLK2_IN                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    GT2_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    ------------------- Receive Ports - Pattern Checker Ports ------------------
    GT2_RXPRBSERR_OUT                       : out  std_logic;
    GT2_RXPRBSSEL_IN                        : in   std_logic_vector(2 downto 0);
    ------------------- Receive Ports - Pattern Checker ports ------------------
    GT2_RXPRBSCNTRESET_IN                   : in   std_logic;
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    GT2_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT2_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GT2_GTHRXN_IN                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    GT2_RXBYTEISALIGNED_OUT                 : out  std_logic;
    GT2_RXCOMMADET_OUT                      : out  std_logic;
    GT2_RXMCOMMAALIGNEN_IN                  : in   std_logic;
    GT2_RXPCOMMAALIGNEN_IN                  : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    GT2_RXOUTCLK_OUT                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GT2_GTRXRESET_IN                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    GT2_RXPOLARITY_IN                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    GT2_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT2_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    GT2_GTHRXP_IN                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    GT2_RXRESETDONE_OUT                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GT2_GTTXRESET_IN                        : in   std_logic;
    GT2_TXUSERRDY_IN                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    GT2_TXUSRCLK_IN                         : in   std_logic;
    GT2_TXUSRCLK2_IN                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GT2_TXDATA_IN                           : in   std_logic_vector(15 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GT2_GTHTXN_OUT                          : out  std_logic;
    GT2_GTHTXP_OUT                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    GT2_TXOUTCLK_OUT                        : out  std_logic;
    GT2_TXOUTCLKFABRIC_OUT                  : out  std_logic;
    GT2_TXOUTCLKPCS_OUT                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    GT2_TXRESETDONE_OUT                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    GT2_TXPOLARITY_IN                       : in   std_logic;
    ------------------ Transmit Ports - pattern Generator Ports ----------------
    GT2_TXPRBSSEL_IN                        : in   std_logic_vector(2 downto 0);
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    GT2_TXCHARISK_IN                        : in   std_logic_vector(1 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT3  (X1Y35)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    GT3_CPLLFBCLKLOST_OUT                   : out  std_logic;
    GT3_CPLLLOCK_OUT                        : out  std_logic;
    GT3_CPLLLOCKDETCLK_IN                   : in   std_logic;
    GT3_CPLLRESET_IN                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    GT3_GTREFCLK0_IN                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    GT3_DRPADDR_IN                          : in   std_logic_vector(8 downto 0);
    GT3_DRPCLK_IN                           : in   std_logic;
    GT3_DRPDI_IN                            : in   std_logic_vector(15 downto 0);
    GT3_DRPDO_OUT                           : out  std_logic_vector(15 downto 0);
    GT3_DRPEN_IN                            : in   std_logic;
    GT3_DRPRDY_OUT                          : out  std_logic;
    GT3_DRPWE_IN                            : in   std_logic;
    ------------------------------- Loopback Ports -----------------------------
    GT3_LOOPBACK_IN                         : in   std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    GT3_RXUSERRDY_IN                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    GT3_EYESCANDATAERROR_OUT                : out  std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    GT3_RXCDRLOCK_OUT                       : out  std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    GT3_RXUSRCLK_IN                         : in   std_logic;
    GT3_RXUSRCLK2_IN                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    GT3_RXDATA_OUT                          : out  std_logic_vector(15 downto 0);
    ------------------- Receive Ports - Pattern Checker Ports ------------------
    GT3_RXPRBSERR_OUT                       : out  std_logic;
    GT3_RXPRBSSEL_IN                        : in   std_logic_vector(2 downto 0);
    ------------------- Receive Ports - Pattern Checker ports ------------------
    GT3_RXPRBSCNTRESET_IN                   : in   std_logic;
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    GT3_RXDISPERR_OUT                       : out  std_logic_vector(1 downto 0);
    GT3_RXNOTINTABLE_OUT                    : out  std_logic_vector(1 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    GT3_GTHRXN_IN                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    GT3_RXBYTEISALIGNED_OUT                 : out  std_logic;
    GT3_RXCOMMADET_OUT                      : out  std_logic;
    GT3_RXMCOMMAALIGNEN_IN                  : in   std_logic;
    GT3_RXPCOMMAALIGNEN_IN                  : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    GT3_RXOUTCLK_OUT                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    GT3_GTRXRESET_IN                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    GT3_RXPOLARITY_IN                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    GT3_RXCHARISCOMMA_OUT                   : out  std_logic_vector(1 downto 0);
    GT3_RXCHARISK_OUT                       : out  std_logic_vector(1 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    GT3_GTHRXP_IN                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    GT3_RXRESETDONE_OUT                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    GT3_GTTXRESET_IN                        : in   std_logic;
    GT3_TXUSERRDY_IN                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    GT3_TXUSRCLK_IN                         : in   std_logic;
    GT3_TXUSRCLK2_IN                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    GT3_TXDATA_IN                           : in   std_logic_vector(15 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    GT3_GTHTXN_OUT                          : out  std_logic;
    GT3_GTHTXP_OUT                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    GT3_TXOUTCLK_OUT                        : out  std_logic;
    GT3_TXOUTCLKFABRIC_OUT                  : out  std_logic;
    GT3_TXOUTCLKPCS_OUT                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    GT3_TXRESETDONE_OUT                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    GT3_TXPOLARITY_IN                       : in   std_logic;
    ------------------ Transmit Ports - pattern Generator Ports ----------------
    GT3_TXPRBSSEL_IN                        : in   std_logic_vector(2 downto 0);
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    GT3_TXCHARISK_IN                        : in   std_logic_vector(1 downto 0);
   

    --____________________________COMMON PORTS________________________________
    ---------------------- Common Block  - Ref Clock Ports ---------------------
    GT0_GTREFCLK0_COMMON_IN                 : in   std_logic;
    ------------------------- Common Block - QPLL Ports ------------------------
    GT0_QPLLLOCK_OUT                        : out  std_logic;
    GT0_QPLLLOCKDETCLK_IN                   : in   std_logic;
    GT0_QPLLRESET_IN                        : in   std_logic


);
end component;

component xilinx_gth_16b_5g_cpll_GT_USRCLK_SOURCE 
port
(
    Q7_CLK0_GTREFCLK_PAD_N_IN               : in   std_logic;
    Q7_CLK0_GTREFCLK_PAD_P_IN               : in   std_logic;
    Q7_CLK0_GTREFCLK_OUT                    : out  std_logic;
 
    GT0_TXUSRCLK_OUT             : out std_logic;
    GT0_TXUSRCLK2_OUT            : out std_logic;
    GT0_TXOUTCLK_IN              : in  std_logic;
    GT0_RXUSRCLK_OUT             : out std_logic;
    GT0_RXUSRCLK2_OUT            : out std_logic;
    GT0_RXOUTCLK_IN              : in  std_logic;
 
    GT1_TXUSRCLK_OUT             : out std_logic;
    GT1_TXUSRCLK2_OUT            : out std_logic;
    GT1_TXOUTCLK_IN              : in  std_logic;
    GT1_RXUSRCLK_OUT             : out std_logic;
    GT1_RXUSRCLK2_OUT            : out std_logic;
    GT1_RXOUTCLK_IN              : in  std_logic;
 
    GT2_TXUSRCLK_OUT             : out std_logic;
    GT2_TXUSRCLK2_OUT            : out std_logic;
    GT2_TXOUTCLK_IN              : in  std_logic;
    GT2_RXUSRCLK_OUT             : out std_logic;
    GT2_RXUSRCLK2_OUT            : out std_logic;
    GT2_RXOUTCLK_IN              : in  std_logic;
 
    GT3_TXUSRCLK_OUT             : out std_logic;
    GT3_TXUSRCLK2_OUT            : out std_logic;
    GT3_TXOUTCLK_IN              : in  std_logic;
    GT3_RXUSRCLK_OUT             : out std_logic;
    GT3_RXUSRCLK2_OUT            : out std_logic;
    GT3_RXOUTCLK_IN              : in  std_logic;
    DRPCLK_IN                          : in  std_logic;
    DRPCLK_OUT                         : out std_logic
);
end component;





component xilinx_gth_16b_5g_cpll_GT_FRAME_GEN 
generic
(
     WORDS_IN_BRAM    : integer := 512
);
port
(
    -- User Interface
    TX_DATA_OUT             : out   std_logic_vector(79 downto 0);
    TXCTRL_OUT              : out   std_logic_vector(7 downto 0); 
    -- System Interface
    USER_CLK                : in    std_logic;      
    SYSTEM_RESET            : in    std_logic
); 
end component;

component xilinx_gth_16b_5g_cpll_GT_FRAME_CHECK 
generic
(
    RX_DATA_WIDTH            : integer := 16;
    RXCTRL_WIDTH             : integer := 2; 
    WORDS_IN_BRAM            : integer := 256;
    CHANBOND_SEQ_LEN         : integer := 1;
    COMMA_DOUBLE             : std_logic_vector(15 downto 0) := x"f628";
    START_OF_PACKET_CHAR     : std_logic_vector(15 downto 0) := x"02bc"
);
port
(
    -- User Interface
    RX_DATA_IN               : in  std_logic_vector((RX_DATA_WIDTH-1) downto 0);
    RXCTRL_IN                : in  std_logic_vector((RXCTRL_WIDTH-1) downto 0); 
    RXENMCOMMADET_OUT        : out std_logic;
    RXENPCOMMADET_OUT        : out std_logic;
    RX_ENCHAN_SYNC_OUT       : out std_logic;
    RX_CHANBOND_SEQ_IN       : in  std_logic;

    -- Control Interface
    INC_IN                   : in  std_logic; 
    INC_OUT                  : out std_logic; 
    PATTERN_MATCHB_OUT       : out std_logic;
    RESET_ON_ERROR_IN        : in  std_logic;


    -- Error Monitoring
    ERROR_COUNT_OUT          : out std_logic_vector(7 downto 0);

    -- Track Data
    TRACK_DATA_OUT           : out std_logic;

 

    -- System Interface
    USER_CLK                 : in std_logic;       
    SYSTEM_RESET             : in std_logic
);
end component;

-- Chipscope modules
attribute syn_black_box                : boolean;
attribute syn_noprune                  : boolean;


component data_vio
port
(
    control                 : inout std_logic_vector(35 downto 0);
    clk                     : in    std_logic;
    async_in                : in    std_logic_vector(31 downto 0);
    async_out               : out   std_logic_vector(31 downto 0);
    sync_in                 : in    std_logic_vector(31 downto 0);
    sync_out                : out   std_logic_vector(31 downto 0)
);
end component;
attribute syn_black_box of data_vio : component is TRUE;
attribute syn_noprune of data_vio   : component is TRUE;


component icon
port
(
    control0                : inout std_logic_vector(35 downto 0);
    control1                : inout std_logic_vector(35 downto 0);
    control2                : inout std_logic_vector(35 downto 0);
    control3                : inout std_logic_vector(35 downto 0);
    control4                : inout std_logic_vector(35 downto 0);
    control5                : inout std_logic_vector(35 downto 0)
);
end component;
attribute syn_black_box of icon : component is TRUE;
attribute syn_noprune of icon   : component is TRUE;


component ila
port
(
    control                 : inout std_logic_vector(35 downto 0);
    clk                     : in    std_logic;
    trig0                   : in    std_logic_vector(163 downto 0)
);
end component;

--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;

--************************** Register Declarations ****************************

    signal   gt0_txfsmresetdone_i            : std_logic;
    signal   gt0_rxfsmresetdone_i            : std_logic;
    signal   gt0_txfsmresetdone_r            : std_logic;
    signal   gt0_txfsmresetdone_r2           : std_logic;
    signal   gt0_rxresetdone_r               : std_logic;
    signal   gt0_rxresetdone_r2              : std_logic;
    signal   gt0_rxresetdone_r3              : std_logic;


    signal   gt1_txfsmresetdone_i            : std_logic;
    signal   gt1_rxfsmresetdone_i            : std_logic;
    signal   gt1_txfsmresetdone_r            : std_logic;
    signal   gt1_txfsmresetdone_r2           : std_logic;
    signal   gt1_rxresetdone_r               : std_logic;
    signal   gt1_rxresetdone_r2              : std_logic;
    signal   gt1_rxresetdone_r3              : std_logic;


    signal   gt2_txfsmresetdone_i            : std_logic;
    signal   gt2_rxfsmresetdone_i            : std_logic;
    signal   gt2_txfsmresetdone_r            : std_logic;
    signal   gt2_txfsmresetdone_r2           : std_logic;
    signal   gt2_rxresetdone_r               : std_logic;
    signal   gt2_rxresetdone_r2              : std_logic;
    signal   gt2_rxresetdone_r3              : std_logic;


    signal   gt3_txfsmresetdone_i            : std_logic;
    signal   gt3_rxfsmresetdone_i            : std_logic;
    signal   gt3_txfsmresetdone_r            : std_logic;
    signal   gt3_txfsmresetdone_r2           : std_logic;
    signal   gt3_rxresetdone_r               : std_logic;
    signal   gt3_rxresetdone_r2              : std_logic;
    signal   gt3_rxresetdone_r3              : std_logic;



--**************************** Wire Declarations ******************************
    -------------------------- GT Wrapper Wires ------------------------------
    --________________________________________________________________________
    --________________________________________________________________________
    --GT0   (X1Y32)

    --------------------------------- CPLL Ports -------------------------------
    signal  gt0_cpllfbclklost_i             : std_logic;
    signal  gt0_cplllock_i                  : std_logic;
    signal  gt0_cpllrefclklost_i            : std_logic;
    signal  gt0_cpllreset_i                 : std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt0_drpaddr_i                   : std_logic_vector(8 downto 0);
    signal  gt0_drpdi_i                     : std_logic_vector(15 downto 0);
    signal  gt0_drpdo_i                     : std_logic_vector(15 downto 0);
    signal  gt0_drpen_i                     : std_logic;
    signal  gt0_drprdy_i                    : std_logic;
    signal  gt0_drpwe_i                     : std_logic;
    ------------------------------- Loopback Ports -----------------------------
    signal  gt0_loopback_i                  : std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt0_rxuserrdy_i                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt0_eyescandataerror_i          : std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    signal  gt0_rxcdrlock_i                 : std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt0_rxdata_i                    : std_logic_vector(15 downto 0);
    ------------------- Receive Ports - Pattern Checker Ports ------------------
    signal  gt0_rxprbserr_i                 : std_logic;
    signal  gt0_rxprbssel_i                 : std_logic_vector(2 downto 0);
    ------------------- Receive Ports - Pattern Checker ports ------------------
    signal  gt0_rxprbscntreset_i            : std_logic;
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt0_rxdisperr_i                 : std_logic_vector(1 downto 0);
    signal  gt0_rxnotintable_i              : std_logic_vector(1 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt0_gthrxn_i                    : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt0_rxbyteisaligned_i           : std_logic;
    signal  gt0_rxcommadet_i                : std_logic;
    signal  gt0_rxmcommaalignen_i           : std_logic;
    signal  gt0_rxpcommaalignen_i           : std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt0_rxoutclk_i                  : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt0_gtrxreset_i                 : std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    signal  gt0_rxpolarity_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt0_rxchariscomma_i             : std_logic_vector(1 downto 0);
    signal  gt0_rxcharisk_i                 : std_logic_vector(1 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt0_gthrxp_i                    : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt0_rxresetdone_i               : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt0_gttxreset_i                 : std_logic;
    signal  gt0_txuserrdy_i                 : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt0_txdata_i                    : std_logic_vector(15 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt0_gthtxn_i                    : std_logic;
    signal  gt0_gthtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt0_txoutclk_i                  : std_logic;
    signal  gt0_txoutclkfabric_i            : std_logic;
    signal  gt0_txoutclkpcs_i               : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt0_txresetdone_i               : std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    signal  gt0_txpolarity_i                : std_logic;
    ------------------ Transmit Ports - pattern Generator Ports ----------------
    signal  gt0_txprbssel_i                 : std_logic_vector(2 downto 0);
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt0_txcharisk_i                 : std_logic_vector(1 downto 0);


    --________________________________________________________________________
    --________________________________________________________________________
    --GT1   (X1Y33)

    --------------------------------- CPLL Ports -------------------------------
    signal  gt1_cpllfbclklost_i             : std_logic;
    signal  gt1_cplllock_i                  : std_logic;
    signal  gt1_cpllrefclklost_i            : std_logic;
    signal  gt1_cpllreset_i                 : std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt1_drpaddr_i                   : std_logic_vector(8 downto 0);
    signal  gt1_drpdi_i                     : std_logic_vector(15 downto 0);
    signal  gt1_drpdo_i                     : std_logic_vector(15 downto 0);
    signal  gt1_drpen_i                     : std_logic;
    signal  gt1_drprdy_i                    : std_logic;
    signal  gt1_drpwe_i                     : std_logic;
    ------------------------------- Loopback Ports -----------------------------
    signal  gt1_loopback_i                  : std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt1_rxuserrdy_i                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt1_eyescandataerror_i          : std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    signal  gt1_rxcdrlock_i                 : std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt1_rxdata_i                    : std_logic_vector(15 downto 0);
    ------------------- Receive Ports - Pattern Checker Ports ------------------
    signal  gt1_rxprbserr_i                 : std_logic;
    signal  gt1_rxprbssel_i                 : std_logic_vector(2 downto 0);
    ------------------- Receive Ports - Pattern Checker ports ------------------
    signal  gt1_rxprbscntreset_i            : std_logic;
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt1_rxdisperr_i                 : std_logic_vector(1 downto 0);
    signal  gt1_rxnotintable_i              : std_logic_vector(1 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt1_gthrxn_i                    : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt1_rxbyteisaligned_i           : std_logic;
    signal  gt1_rxcommadet_i                : std_logic;
    signal  gt1_rxmcommaalignen_i           : std_logic;
    signal  gt1_rxpcommaalignen_i           : std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt1_rxoutclk_i                  : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt1_gtrxreset_i                 : std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    signal  gt1_rxpolarity_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt1_rxchariscomma_i             : std_logic_vector(1 downto 0);
    signal  gt1_rxcharisk_i                 : std_logic_vector(1 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt1_gthrxp_i                    : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt1_rxresetdone_i               : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt1_gttxreset_i                 : std_logic;
    signal  gt1_txuserrdy_i                 : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt1_txdata_i                    : std_logic_vector(15 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt1_gthtxn_i                    : std_logic;
    signal  gt1_gthtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt1_txoutclk_i                  : std_logic;
    signal  gt1_txoutclkfabric_i            : std_logic;
    signal  gt1_txoutclkpcs_i               : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt1_txresetdone_i               : std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    signal  gt1_txpolarity_i                : std_logic;
    ------------------ Transmit Ports - pattern Generator Ports ----------------
    signal  gt1_txprbssel_i                 : std_logic_vector(2 downto 0);
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt1_txcharisk_i                 : std_logic_vector(1 downto 0);


    --________________________________________________________________________
    --________________________________________________________________________
    --GT2   (X1Y34)

    --------------------------------- CPLL Ports -------------------------------
    signal  gt2_cpllfbclklost_i             : std_logic;
    signal  gt2_cplllock_i                  : std_logic;
    signal  gt2_cpllrefclklost_i            : std_logic;
    signal  gt2_cpllreset_i                 : std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt2_drpaddr_i                   : std_logic_vector(8 downto 0);
    signal  gt2_drpdi_i                     : std_logic_vector(15 downto 0);
    signal  gt2_drpdo_i                     : std_logic_vector(15 downto 0);
    signal  gt2_drpen_i                     : std_logic;
    signal  gt2_drprdy_i                    : std_logic;
    signal  gt2_drpwe_i                     : std_logic;
    ------------------------------- Loopback Ports -----------------------------
    signal  gt2_loopback_i                  : std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt2_rxuserrdy_i                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt2_eyescandataerror_i          : std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    signal  gt2_rxcdrlock_i                 : std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt2_rxdata_i                    : std_logic_vector(15 downto 0);
    ------------------- Receive Ports - Pattern Checker Ports ------------------
    signal  gt2_rxprbserr_i                 : std_logic;
    signal  gt2_rxprbssel_i                 : std_logic_vector(2 downto 0);
    ------------------- Receive Ports - Pattern Checker ports ------------------
    signal  gt2_rxprbscntreset_i            : std_logic;
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt2_rxdisperr_i                 : std_logic_vector(1 downto 0);
    signal  gt2_rxnotintable_i              : std_logic_vector(1 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt2_gthrxn_i                    : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt2_rxbyteisaligned_i           : std_logic;
    signal  gt2_rxcommadet_i                : std_logic;
    signal  gt2_rxmcommaalignen_i           : std_logic;
    signal  gt2_rxpcommaalignen_i           : std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt2_rxoutclk_i                  : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt2_gtrxreset_i                 : std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    signal  gt2_rxpolarity_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt2_rxchariscomma_i             : std_logic_vector(1 downto 0);
    signal  gt2_rxcharisk_i                 : std_logic_vector(1 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt2_gthrxp_i                    : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt2_rxresetdone_i               : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt2_gttxreset_i                 : std_logic;
    signal  gt2_txuserrdy_i                 : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt2_txdata_i                    : std_logic_vector(15 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt2_gthtxn_i                    : std_logic;
    signal  gt2_gthtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt2_txoutclk_i                  : std_logic;
    signal  gt2_txoutclkfabric_i            : std_logic;
    signal  gt2_txoutclkpcs_i               : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt2_txresetdone_i               : std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    signal  gt2_txpolarity_i                : std_logic;
    ------------------ Transmit Ports - pattern Generator Ports ----------------
    signal  gt2_txprbssel_i                 : std_logic_vector(2 downto 0);
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt2_txcharisk_i                 : std_logic_vector(1 downto 0);


    --________________________________________________________________________
    --________________________________________________________________________
    --GT3   (X1Y35)

    --------------------------------- CPLL Ports -------------------------------
    signal  gt3_cpllfbclklost_i             : std_logic;
    signal  gt3_cplllock_i                  : std_logic;
    signal  gt3_cpllrefclklost_i            : std_logic;
    signal  gt3_cpllreset_i                 : std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt3_drpaddr_i                   : std_logic_vector(8 downto 0);
    signal  gt3_drpdi_i                     : std_logic_vector(15 downto 0);
    signal  gt3_drpdo_i                     : std_logic_vector(15 downto 0);
    signal  gt3_drpen_i                     : std_logic;
    signal  gt3_drprdy_i                    : std_logic;
    signal  gt3_drpwe_i                     : std_logic;
    ------------------------------- Loopback Ports -----------------------------
    signal  gt3_loopback_i                  : std_logic_vector(2 downto 0);
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt3_rxuserrdy_i                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt3_eyescandataerror_i          : std_logic;
    ------------------------- Receive Ports - CDR Ports ------------------------
    signal  gt3_rxcdrlock_i                 : std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    signal  gt3_rxdata_i                    : std_logic_vector(15 downto 0);
    ------------------- Receive Ports - Pattern Checker Ports ------------------
    signal  gt3_rxprbserr_i                 : std_logic;
    signal  gt3_rxprbssel_i                 : std_logic_vector(2 downto 0);
    ------------------- Receive Ports - Pattern Checker ports ------------------
    signal  gt3_rxprbscntreset_i            : std_logic;
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt3_rxdisperr_i                 : std_logic_vector(1 downto 0);
    signal  gt3_rxnotintable_i              : std_logic_vector(1 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt3_gthrxn_i                    : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt3_rxbyteisaligned_i           : std_logic;
    signal  gt3_rxcommadet_i                : std_logic;
    signal  gt3_rxmcommaalignen_i           : std_logic;
    signal  gt3_rxpcommaalignen_i           : std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt3_rxoutclk_i                  : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt3_gtrxreset_i                 : std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    signal  gt3_rxpolarity_i                : std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    signal  gt3_rxchariscomma_i             : std_logic_vector(1 downto 0);
    signal  gt3_rxcharisk_i                 : std_logic_vector(1 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    signal  gt3_gthrxp_i                    : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt3_rxresetdone_i               : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt3_gttxreset_i                 : std_logic;
    signal  gt3_txuserrdy_i                 : std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  gt3_txdata_i                    : std_logic_vector(15 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    signal  gt3_gthtxn_i                    : std_logic;
    signal  gt3_gthtxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt3_txoutclk_i                  : std_logic;
    signal  gt3_txoutclkfabric_i            : std_logic;
    signal  gt3_txoutclkpcs_i               : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt3_txresetdone_i               : std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    signal  gt3_txpolarity_i                : std_logic;
    ------------------ Transmit Ports - pattern Generator Ports ----------------
    signal  gt3_txprbssel_i                 : std_logic_vector(2 downto 0);
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    signal  gt3_txcharisk_i                 : std_logic_vector(1 downto 0);



    --____________________________COMMON PORTS________________________________
    ------------------------- Common Block - QPLL Ports ------------------------
    signal  gt0_qplllock_i                  : std_logic;
    signal  gt0_qpllrefclklost_i            : std_logic;
    signal  gt0_qpllreset_i                 : std_logic;



    ------------------------------- Global Signals -----------------------------
    signal  gt0_tx_system_reset_c           : std_logic;
    signal  gt0_rx_system_reset_c           : std_logic;
    signal  gt1_tx_system_reset_c           : std_logic;
    signal  gt1_rx_system_reset_c           : std_logic;
    signal  gt2_tx_system_reset_c           : std_logic;
    signal  gt2_rx_system_reset_c           : std_logic;
    signal  gt3_tx_system_reset_c           : std_logic;
    signal  gt3_rx_system_reset_c           : std_logic;
    signal  tied_to_ground_i                : std_logic;
    signal  tied_to_ground_vec_i            : std_logic_vector(63 downto 0);
    signal  tied_to_vcc_i                   : std_logic;
    signal  tied_to_vcc_vec_i               : std_logic_vector(7 downto 0);
    signal  drpclk_in_i                     : std_logic;
 
    signal  GTTXRESET_IN                    : std_logic;
    signal  GTRXRESET_IN                    : std_logic;
    signal  CPLLRESET_IN                    : std_logic;
    signal  QPLLRESET_IN                    : std_logic;

   ------------------------------- User Clocks ---------------------------------
    attribute keep: string;
    signal    gt0_txusrclk_i                  : std_logic; 
    signal    gt0_txusrclk2_i                 : std_logic; 
    signal    gt0_rxusrclk_i                  : std_logic; 
    signal    gt0_rxusrclk2_i                 : std_logic; 
    attribute keep of gt0_txusrclk_i : signal is "true";
    attribute keep of gt0_txusrclk2_i : signal is "true";
    attribute keep of gt0_rxusrclk_i : signal is "true";
    attribute keep of gt0_rxusrclk2_i : signal is "true";
    signal    gt1_txusrclk_i                  : std_logic; 
    signal    gt1_txusrclk2_i                 : std_logic; 
    signal    gt1_rxusrclk_i                  : std_logic; 
    signal    gt1_rxusrclk2_i                 : std_logic; 
    attribute keep of gt1_txusrclk_i : signal is "true";
    attribute keep of gt1_txusrclk2_i : signal is "true";
    attribute keep of gt1_rxusrclk_i : signal is "true";
    attribute keep of gt1_rxusrclk2_i : signal is "true";
    signal    gt2_txusrclk_i                  : std_logic; 
    signal    gt2_txusrclk2_i                 : std_logic; 
    signal    gt2_rxusrclk_i                  : std_logic; 
    signal    gt2_rxusrclk2_i                 : std_logic; 
    attribute keep of gt2_txusrclk_i : signal is "true";
    attribute keep of gt2_txusrclk2_i : signal is "true";
    attribute keep of gt2_rxusrclk_i : signal is "true";
    attribute keep of gt2_rxusrclk2_i : signal is "true";
    signal    gt3_txusrclk_i                  : std_logic; 
    signal    gt3_txusrclk2_i                 : std_logic; 
    signal    gt3_rxusrclk_i                  : std_logic; 
    signal    gt3_rxusrclk2_i                 : std_logic; 
    attribute keep of gt3_txusrclk_i : signal is "true";
    attribute keep of gt3_txusrclk2_i : signal is "true";
    attribute keep of gt3_rxusrclk_i : signal is "true";
    attribute keep of gt3_rxusrclk2_i : signal is "true";
 



    ----------------------------- Reference Clocks ----------------------------
    
    signal    q7_clk0_refclk_i                : std_logic;


    ----------------------- Frame check/gen Module Signals --------------------
    
    signal    gt0_matchn_i                    : std_logic;
    
    signal    gt0_txcharisk_float_i           : std_logic_vector(5 downto 0);
    
    signal    gt0_txdata_float16_i            : std_logic_vector(15 downto 0);
    signal    gt0_txdata_float_i              : std_logic_vector(47 downto 0);
    
    signal    gt0_track_data_i                : std_logic;
    signal    gt0_block_sync_i                : std_logic;
    signal    gt0_error_count_i               : std_logic_vector(7 downto 0);
    signal    gt0_frame_check_reset_i         : std_logic;
    signal    gt0_inc_in_i                    : std_logic;
    signal    gt0_inc_out_i                   : std_logic;
    signal    gt0_unscrambled_data_i          : std_logic_vector(15 downto 0);

    signal    gt1_matchn_i                    : std_logic;
    
    signal    gt1_txcharisk_float_i           : std_logic_vector(5 downto 0);
    
    signal    gt1_txdata_float16_i            : std_logic_vector(15 downto 0);
    signal    gt1_txdata_float_i              : std_logic_vector(47 downto 0);
    
    signal    gt1_track_data_i                : std_logic;
    signal    gt1_block_sync_i                : std_logic;
    signal    gt1_error_count_i               : std_logic_vector(7 downto 0);
    signal    gt1_frame_check_reset_i         : std_logic;
    signal    gt1_inc_in_i                    : std_logic;
    signal    gt1_inc_out_i                   : std_logic;
    signal    gt1_unscrambled_data_i          : std_logic_vector(15 downto 0);

    signal    gt2_matchn_i                    : std_logic;
    
    signal    gt2_txcharisk_float_i           : std_logic_vector(5 downto 0);
    
    signal    gt2_txdata_float16_i            : std_logic_vector(15 downto 0);
    signal    gt2_txdata_float_i              : std_logic_vector(47 downto 0);
    
    signal    gt2_track_data_i                : std_logic;
    signal    gt2_block_sync_i                : std_logic;
    signal    gt2_error_count_i               : std_logic_vector(7 downto 0);
    signal    gt2_frame_check_reset_i         : std_logic;
    signal    gt2_inc_in_i                    : std_logic;
    signal    gt2_inc_out_i                   : std_logic;
    signal    gt2_unscrambled_data_i          : std_logic_vector(15 downto 0);

    signal    gt3_matchn_i                    : std_logic;
    
    signal    gt3_txcharisk_float_i           : std_logic_vector(5 downto 0);
    
    signal    gt3_txdata_float16_i            : std_logic_vector(15 downto 0);
    signal    gt3_txdata_float_i              : std_logic_vector(47 downto 0);
    
    signal    gt3_track_data_i                : std_logic;
    signal    gt3_block_sync_i                : std_logic;
    signal    gt3_error_count_i               : std_logic_vector(7 downto 0);
    signal    gt3_frame_check_reset_i         : std_logic;
    signal    gt3_inc_in_i                    : std_logic;
    signal    gt3_inc_out_i                   : std_logic;
    signal    gt3_unscrambled_data_i          : std_logic_vector(15 downto 0);

    signal    reset_on_data_error_i           : std_logic;
    signal    track_data_out_i                : std_logic;
   

    ----------------------- Chipscope Signals ---------------------------------

    signal  tx_data_vio_control_i           : std_logic_vector(35 downto 0);
    signal  rx_data_vio_control_i           : std_logic_vector(35 downto 0);
    signal  shared_vio_control_i            : std_logic_vector(35 downto 0);
    signal  ila_control_i                   : std_logic_vector(35 downto 0);
    signal  channel_drp_vio_control_i       : std_logic_vector(35 downto 0);
    signal  common_drp_vio_control_i        : std_logic_vector(35 downto 0);
    signal  tx_data_vio_async_in_i          : std_logic_vector(31 downto 0);
    signal  tx_data_vio_sync_in_i           : std_logic_vector(31 downto 0);
    signal  tx_data_vio_async_out_i         : std_logic_vector(31 downto 0);
    signal  tx_data_vio_sync_out_i          : std_logic_vector(31 downto 0);
    signal  rx_data_vio_async_in_i          : std_logic_vector(31 downto 0);
    signal  rx_data_vio_sync_in_i           : std_logic_vector(31 downto 0);
    signal  rx_data_vio_async_out_i         : std_logic_vector(31 downto 0);
    signal  rx_data_vio_sync_out_i          : std_logic_vector(31 downto 0);
    signal  shared_vio_in_i                 : std_logic_vector(31 downto 0);
    signal  shared_vio_out_i                : std_logic_vector(31 downto 0);
    signal  ila_in_i                        : std_logic_vector(163 downto 0);
    signal  channel_drp_vio_async_in_i      : std_logic_vector(31 downto 0);
    signal  channel_drp_vio_sync_in_i       : std_logic_vector(31 downto 0);
    signal  channel_drp_vio_async_out_i     : std_logic_vector(31 downto 0);
    signal  channel_drp_vio_sync_out_i      : std_logic_vector(31 downto 0);
    signal  common_drp_vio_async_in_i       : std_logic_vector(31 downto 0);
    signal  common_drp_vio_sync_in_i        : std_logic_vector(31 downto 0);
    signal  common_drp_vio_async_out_i      : std_logic_vector(31 downto 0);
    signal  common_drp_vio_sync_out_i       : std_logic_vector(31 downto 0);

    signal  gt0_tx_data_vio_async_in_i      : std_logic_vector(31 downto 0);
    signal  gt0_tx_data_vio_sync_in_i       : std_logic_vector(31 downto 0);
    signal  gt0_tx_data_vio_async_out_i     : std_logic_vector(31 downto 0);
    signal  gt0_tx_data_vio_sync_out_i      : std_logic_vector(31 downto 0);
    signal  gt0_rx_data_vio_async_in_i      : std_logic_vector(31 downto 0);
    signal  gt0_rx_data_vio_sync_in_i       : std_logic_vector(31 downto 0);
    signal  gt0_rx_data_vio_async_out_i     : std_logic_vector(31 downto 0);
    signal  gt0_rx_data_vio_sync_out_i      : std_logic_vector(31 downto 0);
    signal  gt0_ila_in_i                    : std_logic_vector(163 downto 0);
    signal  gt0_channel_drp_vio_async_in_i  : std_logic_vector(31 downto 0);
    signal  gt0_channel_drp_vio_sync_in_i   : std_logic_vector(31 downto 0);
    signal  gt0_channel_drp_vio_async_out_i : std_logic_vector(31 downto 0);
    signal  gt0_channel_drp_vio_sync_out_i  : std_logic_vector(31 downto 0);
    signal  gt0_common_drp_vio_async_in_i   : std_logic_vector(31 downto 0);
    signal  gt0_common_drp_vio_sync_in_i    : std_logic_vector(31 downto 0);
    signal  gt0_common_drp_vio_async_out_i  : std_logic_vector(31 downto 0);
    signal  gt0_common_drp_vio_sync_out_i   : std_logic_vector(31 downto 0);

    signal  gt1_tx_data_vio_async_in_i      : std_logic_vector(31 downto 0);
    signal  gt1_tx_data_vio_sync_in_i       : std_logic_vector(31 downto 0);
    signal  gt1_tx_data_vio_async_out_i     : std_logic_vector(31 downto 0);
    signal  gt1_tx_data_vio_sync_out_i      : std_logic_vector(31 downto 0);
    signal  gt1_rx_data_vio_async_in_i      : std_logic_vector(31 downto 0);
    signal  gt1_rx_data_vio_sync_in_i       : std_logic_vector(31 downto 0);
    signal  gt1_rx_data_vio_async_out_i     : std_logic_vector(31 downto 0);
    signal  gt1_rx_data_vio_sync_out_i      : std_logic_vector(31 downto 0);
    signal  gt1_ila_in_i                    : std_logic_vector(163 downto 0);
    signal  gt1_channel_drp_vio_async_in_i  : std_logic_vector(31 downto 0);
    signal  gt1_channel_drp_vio_sync_in_i   : std_logic_vector(31 downto 0);
    signal  gt1_channel_drp_vio_async_out_i : std_logic_vector(31 downto 0);
    signal  gt1_channel_drp_vio_sync_out_i  : std_logic_vector(31 downto 0);
    signal  gt1_common_drp_vio_async_in_i   : std_logic_vector(31 downto 0);
    signal  gt1_common_drp_vio_sync_in_i    : std_logic_vector(31 downto 0);
    signal  gt1_common_drp_vio_async_out_i  : std_logic_vector(31 downto 0);
    signal  gt1_common_drp_vio_sync_out_i   : std_logic_vector(31 downto 0);

    signal  gt2_tx_data_vio_async_in_i      : std_logic_vector(31 downto 0);
    signal  gt2_tx_data_vio_sync_in_i       : std_logic_vector(31 downto 0);
    signal  gt2_tx_data_vio_async_out_i     : std_logic_vector(31 downto 0);
    signal  gt2_tx_data_vio_sync_out_i      : std_logic_vector(31 downto 0);
    signal  gt2_rx_data_vio_async_in_i      : std_logic_vector(31 downto 0);
    signal  gt2_rx_data_vio_sync_in_i       : std_logic_vector(31 downto 0);
    signal  gt2_rx_data_vio_async_out_i     : std_logic_vector(31 downto 0);
    signal  gt2_rx_data_vio_sync_out_i      : std_logic_vector(31 downto 0);
    signal  gt2_ila_in_i                    : std_logic_vector(163 downto 0);
    signal  gt2_channel_drp_vio_async_in_i  : std_logic_vector(31 downto 0);
    signal  gt2_channel_drp_vio_sync_in_i   : std_logic_vector(31 downto 0);
    signal  gt2_channel_drp_vio_async_out_i : std_logic_vector(31 downto 0);
    signal  gt2_channel_drp_vio_sync_out_i  : std_logic_vector(31 downto 0);
    signal  gt2_common_drp_vio_async_in_i   : std_logic_vector(31 downto 0);
    signal  gt2_common_drp_vio_sync_in_i    : std_logic_vector(31 downto 0);
    signal  gt2_common_drp_vio_async_out_i  : std_logic_vector(31 downto 0);
    signal  gt2_common_drp_vio_sync_out_i   : std_logic_vector(31 downto 0);

    signal  gt3_tx_data_vio_async_in_i      : std_logic_vector(31 downto 0);
    signal  gt3_tx_data_vio_sync_in_i       : std_logic_vector(31 downto 0);
    signal  gt3_tx_data_vio_async_out_i     : std_logic_vector(31 downto 0);
    signal  gt3_tx_data_vio_sync_out_i      : std_logic_vector(31 downto 0);
    signal  gt3_rx_data_vio_async_in_i      : std_logic_vector(31 downto 0);
    signal  gt3_rx_data_vio_sync_in_i       : std_logic_vector(31 downto 0);
    signal  gt3_rx_data_vio_async_out_i     : std_logic_vector(31 downto 0);
    signal  gt3_rx_data_vio_sync_out_i      : std_logic_vector(31 downto 0);
    signal  gt3_ila_in_i                    : std_logic_vector(163 downto 0);
    signal  gt3_channel_drp_vio_async_in_i  : std_logic_vector(31 downto 0);
    signal  gt3_channel_drp_vio_sync_in_i   : std_logic_vector(31 downto 0);
    signal  gt3_channel_drp_vio_async_out_i : std_logic_vector(31 downto 0);
    signal  gt3_channel_drp_vio_sync_out_i  : std_logic_vector(31 downto 0);
    signal  gt3_common_drp_vio_async_in_i   : std_logic_vector(31 downto 0);
    signal  gt3_common_drp_vio_sync_in_i    : std_logic_vector(31 downto 0);
    signal  gt3_common_drp_vio_async_out_i  : std_logic_vector(31 downto 0);
    signal  gt3_common_drp_vio_sync_out_i   : std_logic_vector(31 downto 0);


    signal    gttxreset_i                     : std_logic;
    signal    gtrxreset_i                     : std_logic;
    signal    mux_sel_i                       : std_logic_vector(1 downto 0);

    signal    user_tx_reset_i                 : std_logic;
    signal    user_rx_reset_i                 : std_logic;
    signal    tx_vio_clk_i                    : std_logic;
    signal    tx_vio_clk_mux_out_i            : std_logic;    
    signal    rx_vio_ila_clk_i                : std_logic;
    signal    rx_vio_ila_clk_mux_out_i        : std_logic;    

    
    signal    cpllreset_i                     : std_logic;
    


   function and_reduce(arg: std_logic_vector) return std_logic is
   variable result: std_logic;
    begin
   result := '1';
   for i in arg'range loop
       result := result and arg(i);
   end loop;
        return result;
    end;


--**************************** Main Body of Code *******************************
begin

    --  Static signal Assigments
    tied_to_ground_i                             <= '0';
    tied_to_ground_vec_i                         <= x"0000000000000000";
    tied_to_vcc_i                                <= '1';
    tied_to_vcc_vec_i                            <= x"ff";

    
  
    
  
    
  
    
  

    gt0_usrclk_source : xilinx_gth_16b_5g_cpll_GT_USRCLK_SOURCE
    port map
    (
        Q7_CLK0_GTREFCLK_PAD_N_IN       =>      Q7_CLK0_GTREFCLK_PAD_N_IN,
        Q7_CLK0_GTREFCLK_PAD_P_IN       =>      Q7_CLK0_GTREFCLK_PAD_P_IN,
        Q7_CLK0_GTREFCLK_OUT            =>      q7_clk0_refclk_i,
 
        GT0_TXUSRCLK_OUT                =>      gt0_txusrclk_i,
        GT0_TXUSRCLK2_OUT               =>      gt0_txusrclk2_i,
        GT0_TXOUTCLK_IN                 =>      gt0_txoutclk_i,
        GT0_RXUSRCLK_OUT                =>      gt0_rxusrclk_i,
        GT0_RXUSRCLK2_OUT               =>      gt0_rxusrclk2_i,
        GT0_RXOUTCLK_IN                 =>      gt0_rxoutclk_i,
 
        GT1_TXUSRCLK_OUT                =>      gt1_txusrclk_i,
        GT1_TXUSRCLK2_OUT               =>      gt1_txusrclk2_i,
        GT1_TXOUTCLK_IN                 =>      gt1_txoutclk_i,
        GT1_RXUSRCLK_OUT                =>      gt1_rxusrclk_i,
        GT1_RXUSRCLK2_OUT               =>      gt1_rxusrclk2_i,
        GT1_RXOUTCLK_IN                 =>      gt1_rxoutclk_i,
 
        GT2_TXUSRCLK_OUT                =>      gt2_txusrclk_i,
        GT2_TXUSRCLK2_OUT               =>      gt2_txusrclk2_i,
        GT2_TXOUTCLK_IN                 =>      gt2_txoutclk_i,
        GT2_RXUSRCLK_OUT                =>      gt2_rxusrclk_i,
        GT2_RXUSRCLK2_OUT               =>      gt2_rxusrclk2_i,
        GT2_RXOUTCLK_IN                 =>      gt2_rxoutclk_i,
 
        GT3_TXUSRCLK_OUT                =>      gt3_txusrclk_i,
        GT3_TXUSRCLK2_OUT               =>      gt3_txusrclk2_i,
        GT3_TXOUTCLK_IN                 =>      gt3_txoutclk_i,
        GT3_RXUSRCLK_OUT                =>      gt3_rxusrclk_i,
        GT3_RXUSRCLK2_OUT               =>      gt3_rxusrclk2_i,
        GT3_RXOUTCLK_IN                 =>      gt3_rxoutclk_i,
        DRPCLK_IN                       =>      DRP_CLK_IN,
        DRPCLK_OUT                      =>      drpclk_in_i

    );


    ----------------------------- The GT Wrapper -----------------------------
    
    -- Use the instantiation template in the example directory to add the GT wrapper to your design.
    -- In this example, the wrapper is wired up for basic operation with a frame generator and frame 
    -- checker. The GTs will reset, then attempt to align and transmit data. If channel bonding is 
    -- enabled, bonding should occur after alignment.


    xilinx_gth_16b_5g_cpll_init_i : xilinx_gth_16b_5g_cpll_init
    generic map
    (
        EXAMPLE_SIM_GTRESET_SPEEDUP     =>      EXAMPLE_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION              =>      EXAMPLE_SIMULATION,
        STABLE_CLOCK_PERIOD             =>      STABLE_CLOCK_PERIOD,
        EXAMPLE_USE_CHIPSCOPE           =>      EXAMPLE_USE_CHIPSCOPE
    )
    port map
    (
        SYSCLK_IN                       =>      drpclk_in_i,
        SOFT_RESET_IN                   =>      tied_to_ground_i,
        DONT_RESET_ON_DATA_ERROR_IN     =>      tied_to_ground_i,
        GT0_TX_FSM_RESET_DONE_OUT       =>      gt0_txfsmresetdone_i,
        GT0_RX_FSM_RESET_DONE_OUT       =>      gt0_rxfsmresetdone_i,
        GT0_DATA_VALID_IN               =>      gt0_track_data_i,
        GT1_TX_FSM_RESET_DONE_OUT       =>      gt1_txfsmresetdone_i,
        GT1_RX_FSM_RESET_DONE_OUT       =>      gt1_rxfsmresetdone_i,
        GT1_DATA_VALID_IN               =>      gt1_track_data_i,
        GT2_TX_FSM_RESET_DONE_OUT       =>      gt2_txfsmresetdone_i,
        GT2_RX_FSM_RESET_DONE_OUT       =>      gt2_rxfsmresetdone_i,
        GT2_DATA_VALID_IN               =>      gt2_track_data_i,
        GT3_TX_FSM_RESET_DONE_OUT       =>      gt3_txfsmresetdone_i,
        GT3_RX_FSM_RESET_DONE_OUT       =>      gt3_rxfsmresetdone_i,
        GT3_DATA_VALID_IN               =>      gt3_track_data_i,
  
 
 
 

        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT0  (X1Y32)

        --------------------------------- CPLL Ports -------------------------------
        GT0_CPLLFBCLKLOST_OUT           =>      gt0_cpllfbclklost_i,
        GT0_CPLLLOCK_OUT                =>      gt0_cplllock_i,
        GT0_CPLLLOCKDETCLK_IN           =>      drpclk_in_i,
        GT0_CPLLRESET_IN                =>      gt0_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        GT0_GTREFCLK0_IN                =>      q7_clk0_refclk_i,
        ---------------------------- Channel - DRP Ports  --------------------------
        GT0_DRPADDR_IN                  =>      gt0_drpaddr_i,
        GT0_DRPCLK_IN                   =>      drpclk_in_i,
        GT0_DRPDI_IN                    =>      gt0_drpdi_i,
        GT0_DRPDO_OUT                   =>      gt0_drpdo_i,
        GT0_DRPEN_IN                    =>      gt0_drpen_i,
        GT0_DRPRDY_OUT                  =>      gt0_drprdy_i,
        GT0_DRPWE_IN                    =>      gt0_drpwe_i,
        ------------------------------- Loopback Ports -----------------------------
        GT0_LOOPBACK_IN                 =>      "000",
        --------------------- RX Initialization and Reset Ports --------------------
        GT0_RXUSERRDY_IN                =>      gt0_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        GT0_EYESCANDATAERROR_OUT        =>      gt0_eyescandataerror_i,
        ------------------------- Receive Ports - CDR Ports ------------------------
        GT0_RXCDRLOCK_OUT               =>      gt0_rxcdrlock_i,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        GT0_RXUSRCLK_IN                 =>      gt0_rxusrclk_i,
        GT0_RXUSRCLK2_IN                =>      gt0_rxusrclk_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        GT0_RXDATA_OUT                  =>      gt0_rxdata_i,
        ------------------- Receive Ports - Pattern Checker Ports ------------------
        GT0_RXPRBSERR_OUT               =>      gt0_rxprbserr_i,
        GT0_RXPRBSSEL_IN                =>      gt0_rxprbssel_i,
        ------------------- Receive Ports - Pattern Checker ports ------------------
        GT0_RXPRBSCNTRESET_IN           =>      gt0_rxprbscntreset_i,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        GT0_RXDISPERR_OUT               =>      gt0_rxdisperr_i,
        GT0_RXNOTINTABLE_OUT            =>      gt0_rxnotintable_i,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        GT0_GTHRXN_IN                   =>      RXN_IN(0),
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        GT0_RXBYTEISALIGNED_OUT         =>      gt0_rxbyteisaligned_i,
        GT0_RXCOMMADET_OUT              =>      gt0_rxcommadet_i,
        GT0_RXMCOMMAALIGNEN_IN          =>      gt0_rxmcommaalignen_i,
        GT0_RXPCOMMAALIGNEN_IN          =>      gt0_rxpcommaalignen_i,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        GT0_RXOUTCLK_OUT                =>      gt0_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        GT0_GTRXRESET_IN                =>      gt0_gtrxreset_i,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        GT0_RXPOLARITY_IN               =>      gt0_rxpolarity_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        GT0_RXCHARISCOMMA_OUT           =>      gt0_rxchariscomma_i,
        GT0_RXCHARISK_OUT               =>      gt0_rxcharisk_i,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        GT0_GTHRXP_IN                   =>      RXP_IN(0),
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        GT0_RXRESETDONE_OUT             =>      gt0_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        GT0_GTTXRESET_IN                =>      gt0_gttxreset_i,
        GT0_TXUSERRDY_IN                =>      gt0_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        GT0_TXUSRCLK_IN                 =>      gt0_txusrclk_i,
        GT0_TXUSRCLK2_IN                =>      gt0_txusrclk_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        GT0_TXDATA_IN                   =>      gt0_txdata_i,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        GT0_GTHTXN_OUT                  =>      TXN_OUT(0),
        GT0_GTHTXP_OUT                  =>      TXP_OUT(0),
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        GT0_TXOUTCLK_OUT                =>      gt0_txoutclk_i,
        GT0_TXOUTCLKFABRIC_OUT          =>      gt0_txoutclkfabric_i,
        GT0_TXOUTCLKPCS_OUT             =>      gt0_txoutclkpcs_i,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        GT0_TXRESETDONE_OUT             =>      gt0_txresetdone_i,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        GT0_TXPOLARITY_IN               =>      gt0_txpolarity_i,
        ------------------ Transmit Ports - pattern Generator Ports ----------------
        GT0_TXPRBSSEL_IN                =>      gt0_txprbssel_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        GT0_TXCHARISK_IN                =>      gt0_txcharisk_i,


  
 
 
 

        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT1  (X1Y33)

        --------------------------------- CPLL Ports -------------------------------
        GT1_CPLLFBCLKLOST_OUT           =>      gt1_cpllfbclklost_i,
        GT1_CPLLLOCK_OUT                =>      gt1_cplllock_i,
        GT1_CPLLLOCKDETCLK_IN           =>      drpclk_in_i,
        GT1_CPLLRESET_IN                =>      gt1_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        GT1_GTREFCLK0_IN                =>      q7_clk0_refclk_i,
        ---------------------------- Channel - DRP Ports  --------------------------
        GT1_DRPADDR_IN                  =>      gt1_drpaddr_i,
        GT1_DRPCLK_IN                   =>      drpclk_in_i,
        GT1_DRPDI_IN                    =>      gt1_drpdi_i,
        GT1_DRPDO_OUT                   =>      gt1_drpdo_i,
        GT1_DRPEN_IN                    =>      gt1_drpen_i,
        GT1_DRPRDY_OUT                  =>      gt1_drprdy_i,
        GT1_DRPWE_IN                    =>      gt1_drpwe_i,
        ------------------------------- Loopback Ports -----------------------------
        GT1_LOOPBACK_IN                 =>      "000",
        --------------------- RX Initialization and Reset Ports --------------------
        GT1_RXUSERRDY_IN                =>      gt1_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        GT1_EYESCANDATAERROR_OUT        =>      gt1_eyescandataerror_i,
        ------------------------- Receive Ports - CDR Ports ------------------------
        GT1_RXCDRLOCK_OUT               =>      gt1_rxcdrlock_i,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        GT1_RXUSRCLK_IN                 =>      gt1_rxusrclk_i,
        GT1_RXUSRCLK2_IN                =>      gt1_rxusrclk_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        GT1_RXDATA_OUT                  =>      gt1_rxdata_i,
        ------------------- Receive Ports - Pattern Checker Ports ------------------
        GT1_RXPRBSERR_OUT               =>      gt1_rxprbserr_i,
        GT1_RXPRBSSEL_IN                =>      gt1_rxprbssel_i,
        ------------------- Receive Ports - Pattern Checker ports ------------------
        GT1_RXPRBSCNTRESET_IN           =>      gt1_rxprbscntreset_i,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        GT1_RXDISPERR_OUT               =>      gt1_rxdisperr_i,
        GT1_RXNOTINTABLE_OUT            =>      gt1_rxnotintable_i,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        GT1_GTHRXN_IN                   =>      RXN_IN(1),
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        GT1_RXBYTEISALIGNED_OUT         =>      gt1_rxbyteisaligned_i,
        GT1_RXCOMMADET_OUT              =>      gt1_rxcommadet_i,
        GT1_RXMCOMMAALIGNEN_IN          =>      gt1_rxmcommaalignen_i,
        GT1_RXPCOMMAALIGNEN_IN          =>      gt1_rxpcommaalignen_i,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        GT1_RXOUTCLK_OUT                =>      gt1_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        GT1_GTRXRESET_IN                =>      gt1_gtrxreset_i,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        GT1_RXPOLARITY_IN               =>      gt1_rxpolarity_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        GT1_RXCHARISCOMMA_OUT           =>      gt1_rxchariscomma_i,
        GT1_RXCHARISK_OUT               =>      gt1_rxcharisk_i,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        GT1_GTHRXP_IN                   =>      RXP_IN(1),
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        GT1_RXRESETDONE_OUT             =>      gt1_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        GT1_GTTXRESET_IN                =>      gt1_gttxreset_i,
        GT1_TXUSERRDY_IN                =>      gt1_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        GT1_TXUSRCLK_IN                 =>      gt0_txusrclk_i,
        GT1_TXUSRCLK2_IN                =>      gt0_txusrclk_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        GT1_TXDATA_IN                   =>      gt1_txdata_i,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        GT1_GTHTXN_OUT                  =>      TXN_OUT(1),
        GT1_GTHTXP_OUT                  =>      TXP_OUT(1),
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        GT1_TXOUTCLK_OUT                =>      gt1_txoutclk_i,
        GT1_TXOUTCLKFABRIC_OUT          =>      gt1_txoutclkfabric_i,
        GT1_TXOUTCLKPCS_OUT             =>      gt1_txoutclkpcs_i,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        GT1_TXRESETDONE_OUT             =>      gt1_txresetdone_i,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        GT1_TXPOLARITY_IN               =>      gt1_txpolarity_i,
        ------------------ Transmit Ports - pattern Generator Ports ----------------
        GT1_TXPRBSSEL_IN                =>      gt1_txprbssel_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        GT1_TXCHARISK_IN                =>      gt1_txcharisk_i,


  
 
 
 

        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT2  (X1Y34)

        --------------------------------- CPLL Ports -------------------------------
        GT2_CPLLFBCLKLOST_OUT           =>      gt2_cpllfbclklost_i,
        GT2_CPLLLOCK_OUT                =>      gt2_cplllock_i,
        GT2_CPLLLOCKDETCLK_IN           =>      drpclk_in_i,
        GT2_CPLLRESET_IN                =>      gt2_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        GT2_GTREFCLK0_IN                =>      q7_clk0_refclk_i,
        ---------------------------- Channel - DRP Ports  --------------------------
        GT2_DRPADDR_IN                  =>      gt2_drpaddr_i,
        GT2_DRPCLK_IN                   =>      drpclk_in_i,
        GT2_DRPDI_IN                    =>      gt2_drpdi_i,
        GT2_DRPDO_OUT                   =>      gt2_drpdo_i,
        GT2_DRPEN_IN                    =>      gt2_drpen_i,
        GT2_DRPRDY_OUT                  =>      gt2_drprdy_i,
        GT2_DRPWE_IN                    =>      gt2_drpwe_i,
        ------------------------------- Loopback Ports -----------------------------
        GT2_LOOPBACK_IN                 =>      "000",
        --------------------- RX Initialization and Reset Ports --------------------
        GT2_RXUSERRDY_IN                =>      gt2_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        GT2_EYESCANDATAERROR_OUT        =>      gt2_eyescandataerror_i,
        ------------------------- Receive Ports - CDR Ports ------------------------
        GT2_RXCDRLOCK_OUT               =>      gt2_rxcdrlock_i,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        GT2_RXUSRCLK_IN                 =>      gt2_rxusrclk_i,
        GT2_RXUSRCLK2_IN                =>      gt2_rxusrclk_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        GT2_RXDATA_OUT                  =>      gt2_rxdata_i,
        ------------------- Receive Ports - Pattern Checker Ports ------------------
        GT2_RXPRBSERR_OUT               =>      gt2_rxprbserr_i,
        GT2_RXPRBSSEL_IN                =>      gt2_rxprbssel_i,
        ------------------- Receive Ports - Pattern Checker ports ------------------
        GT2_RXPRBSCNTRESET_IN           =>      gt2_rxprbscntreset_i,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        GT2_RXDISPERR_OUT               =>      gt2_rxdisperr_i,
        GT2_RXNOTINTABLE_OUT            =>      gt2_rxnotintable_i,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        GT2_GTHRXN_IN                   =>      RXN_IN(2),
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        GT2_RXBYTEISALIGNED_OUT         =>      gt2_rxbyteisaligned_i,
        GT2_RXCOMMADET_OUT              =>      gt2_rxcommadet_i,
        GT2_RXMCOMMAALIGNEN_IN          =>      gt2_rxmcommaalignen_i,
        GT2_RXPCOMMAALIGNEN_IN          =>      gt2_rxpcommaalignen_i,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        GT2_RXOUTCLK_OUT                =>      gt2_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        GT2_GTRXRESET_IN                =>      gt2_gtrxreset_i,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        GT2_RXPOLARITY_IN               =>      gt2_rxpolarity_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        GT2_RXCHARISCOMMA_OUT           =>      gt2_rxchariscomma_i,
        GT2_RXCHARISK_OUT               =>      gt2_rxcharisk_i,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        GT2_GTHRXP_IN                   =>      RXP_IN(2),
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        GT2_RXRESETDONE_OUT             =>      gt2_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        GT2_GTTXRESET_IN                =>      gt2_gttxreset_i,
        GT2_TXUSERRDY_IN                =>      gt2_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        GT2_TXUSRCLK_IN                 =>      gt0_txusrclk_i,
        GT2_TXUSRCLK2_IN                =>      gt0_txusrclk_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        GT2_TXDATA_IN                   =>      gt2_txdata_i,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        GT2_GTHTXN_OUT                  =>      TXN_OUT(2),
        GT2_GTHTXP_OUT                  =>      TXP_OUT(2),
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        GT2_TXOUTCLK_OUT                =>      gt2_txoutclk_i,
        GT2_TXOUTCLKFABRIC_OUT          =>      gt2_txoutclkfabric_i,
        GT2_TXOUTCLKPCS_OUT             =>      gt2_txoutclkpcs_i,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        GT2_TXRESETDONE_OUT             =>      gt2_txresetdone_i,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        GT2_TXPOLARITY_IN               =>      gt2_txpolarity_i,
        ------------------ Transmit Ports - pattern Generator Ports ----------------
        GT2_TXPRBSSEL_IN                =>      gt2_txprbssel_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        GT2_TXCHARISK_IN                =>      gt2_txcharisk_i,


  
 
 
 

        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT3  (X1Y35)

        --------------------------------- CPLL Ports -------------------------------
        GT3_CPLLFBCLKLOST_OUT           =>      gt3_cpllfbclklost_i,
        GT3_CPLLLOCK_OUT                =>      gt3_cplllock_i,
        GT3_CPLLLOCKDETCLK_IN           =>      drpclk_in_i,
        GT3_CPLLRESET_IN                =>      gt3_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        GT3_GTREFCLK0_IN                =>      q7_clk0_refclk_i,
        ---------------------------- Channel - DRP Ports  --------------------------
        GT3_DRPADDR_IN                  =>      gt3_drpaddr_i,
        GT3_DRPCLK_IN                   =>      drpclk_in_i,
        GT3_DRPDI_IN                    =>      gt3_drpdi_i,
        GT3_DRPDO_OUT                   =>      gt3_drpdo_i,
        GT3_DRPEN_IN                    =>      gt3_drpen_i,
        GT3_DRPRDY_OUT                  =>      gt3_drprdy_i,
        GT3_DRPWE_IN                    =>      gt3_drpwe_i,
        ------------------------------- Loopback Ports -----------------------------
        GT3_LOOPBACK_IN                 =>      "000",
        --------------------- RX Initialization and Reset Ports --------------------
        GT3_RXUSERRDY_IN                =>      gt3_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        GT3_EYESCANDATAERROR_OUT        =>      gt3_eyescandataerror_i,
        ------------------------- Receive Ports - CDR Ports ------------------------
        GT3_RXCDRLOCK_OUT               =>      gt3_rxcdrlock_i,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        GT3_RXUSRCLK_IN                 =>      gt3_rxusrclk_i,
        GT3_RXUSRCLK2_IN                =>      gt3_rxusrclk_i,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        GT3_RXDATA_OUT                  =>      gt3_rxdata_i,
        ------------------- Receive Ports - Pattern Checker Ports ------------------
        GT3_RXPRBSERR_OUT               =>      gt3_rxprbserr_i,
        GT3_RXPRBSSEL_IN                =>      gt3_rxprbssel_i,
        ------------------- Receive Ports - Pattern Checker ports ------------------
        GT3_RXPRBSCNTRESET_IN           =>      gt3_rxprbscntreset_i,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        GT3_RXDISPERR_OUT               =>      gt3_rxdisperr_i,
        GT3_RXNOTINTABLE_OUT            =>      gt3_rxnotintable_i,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        GT3_GTHRXN_IN                   =>      RXN_IN(3),
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        GT3_RXBYTEISALIGNED_OUT         =>      gt3_rxbyteisaligned_i,
        GT3_RXCOMMADET_OUT              =>      gt3_rxcommadet_i,
        GT3_RXMCOMMAALIGNEN_IN          =>      gt3_rxmcommaalignen_i,
        GT3_RXPCOMMAALIGNEN_IN          =>      gt3_rxpcommaalignen_i,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        GT3_RXOUTCLK_OUT                =>      gt3_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        GT3_GTRXRESET_IN                =>      gt3_gtrxreset_i,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        GT3_RXPOLARITY_IN               =>      gt3_rxpolarity_i,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        GT3_RXCHARISCOMMA_OUT           =>      gt3_rxchariscomma_i,
        GT3_RXCHARISK_OUT               =>      gt3_rxcharisk_i,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        GT3_GTHRXP_IN                   =>      RXP_IN(3),
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        GT3_RXRESETDONE_OUT             =>      gt3_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        GT3_GTTXRESET_IN                =>      gt3_gttxreset_i,
        GT3_TXUSERRDY_IN                =>      gt3_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        GT3_TXUSRCLK_IN                 =>      gt0_txusrclk_i,
        GT3_TXUSRCLK2_IN                =>      gt0_txusrclk_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        GT3_TXDATA_IN                   =>      gt3_txdata_i,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        GT3_GTHTXN_OUT                  =>      TXN_OUT(3),
        GT3_GTHTXP_OUT                  =>      TXP_OUT(3),
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        GT3_TXOUTCLK_OUT                =>      gt3_txoutclk_i,
        GT3_TXOUTCLKFABRIC_OUT          =>      gt3_txoutclkfabric_i,
        GT3_TXOUTCLKPCS_OUT             =>      gt3_txoutclkpcs_i,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        GT3_TXRESETDONE_OUT             =>      gt3_txresetdone_i,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        GT3_TXPOLARITY_IN               =>      gt3_txpolarity_i,
        ------------------ Transmit Ports - pattern Generator Ports ----------------
        GT3_TXPRBSSEL_IN                =>      gt3_txprbssel_i,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        GT3_TXCHARISK_IN                =>      gt3_txcharisk_i,




    --____________________________COMMON PORTS________________________________
        ---------------------- Common Block  - Ref Clock Ports ---------------------
        GT0_GTREFCLK0_COMMON_IN         =>      q7_clk0_refclk_i,
        ------------------------- Common Block - QPLL Ports ------------------------
        GT0_QPLLLOCK_OUT                =>      gt0_qplllock_i,
        GT0_QPLLLOCKDETCLK_IN           =>      drpclk_in_i,
        GT0_QPLLRESET_IN                =>      gt0_qpllreset_i

    );


    -------------------------- User Module Resets -----------------------------
    -- All the User Modules i.e. FRAME_GEN, FRAME_CHECK and the sync modules
    -- are held in reset till the RESETDONE goes high. 
    -- The RESETDONE is registered a couple of times on USRCLK2 and connected 
    -- to the reset of the modules
    
    process( gt0_rxusrclk_i,gt0_rxresetdone_i)
    begin
        if(gt0_rxresetdone_i = '0') then
            gt0_rxresetdone_r  <= '0'   after DLY;
            gt0_rxresetdone_r2 <= '0'   after DLY;
        elsif(gt0_rxusrclk_i'event and gt0_rxusrclk_i = '1') then
            gt0_rxresetdone_r  <= gt0_rxresetdone_i   after DLY;
            gt0_rxresetdone_r2 <= gt0_rxresetdone_r   after DLY;
            gt0_rxresetdone_r3  <= gt0_rxresetdone_r2   after DLY;
        end if;
    end process;


    process( gt0_txusrclk_i,gt0_txfsmresetdone_i)
    begin
        if(gt0_txfsmresetdone_i = '0') then
            gt0_txfsmresetdone_r  <= '0'   after DLY;
            gt0_txfsmresetdone_r2 <= '0'   after DLY;
        elsif(gt0_txusrclk_i'event and gt0_txusrclk_i = '1') then
            gt0_txfsmresetdone_r  <= gt0_txfsmresetdone_i   after DLY;
            gt0_txfsmresetdone_r2 <= gt0_txfsmresetdone_r   after DLY;
        end if;
    end process;
    process( gt1_rxusrclk_i,gt1_rxresetdone_i)
    begin
        if(gt1_rxresetdone_i = '0') then
            gt1_rxresetdone_r  <= '0'   after DLY;
            gt1_rxresetdone_r2 <= '0'   after DLY;
        elsif(gt1_rxusrclk_i'event and gt1_rxusrclk_i = '1') then
            gt1_rxresetdone_r  <= gt1_rxresetdone_i   after DLY;
            gt1_rxresetdone_r2 <= gt1_rxresetdone_r   after DLY;
            gt1_rxresetdone_r3  <= gt1_rxresetdone_r2   after DLY;
        end if;
    end process;


    process( gt0_txusrclk_i,gt1_txfsmresetdone_i)
    begin
        if(gt1_txfsmresetdone_i = '0') then
            gt1_txfsmresetdone_r  <= '0'   after DLY;
            gt1_txfsmresetdone_r2 <= '0'   after DLY;
        elsif(gt0_txusrclk_i'event and gt0_txusrclk_i = '1') then
            gt1_txfsmresetdone_r  <= gt1_txfsmresetdone_i   after DLY;
            gt1_txfsmresetdone_r2 <= gt1_txfsmresetdone_r   after DLY;
        end if;
    end process;
    process( gt2_rxusrclk_i,gt2_rxresetdone_i)
    begin
        if(gt2_rxresetdone_i = '0') then
            gt2_rxresetdone_r  <= '0'   after DLY;
            gt2_rxresetdone_r2 <= '0'   after DLY;
        elsif(gt2_rxusrclk_i'event and gt2_rxusrclk_i = '1') then
            gt2_rxresetdone_r  <= gt2_rxresetdone_i   after DLY;
            gt2_rxresetdone_r2 <= gt2_rxresetdone_r   after DLY;
            gt2_rxresetdone_r3  <= gt2_rxresetdone_r2   after DLY;
        end if;
    end process;


    process( gt0_txusrclk_i,gt2_txfsmresetdone_i)
    begin
        if(gt2_txfsmresetdone_i = '0') then
            gt2_txfsmresetdone_r  <= '0'   after DLY;
            gt2_txfsmresetdone_r2 <= '0'   after DLY;
        elsif(gt0_txusrclk_i'event and gt0_txusrclk_i = '1') then
            gt2_txfsmresetdone_r  <= gt2_txfsmresetdone_i   after DLY;
            gt2_txfsmresetdone_r2 <= gt2_txfsmresetdone_r   after DLY;
        end if;
    end process;
    process( gt3_rxusrclk_i,gt3_rxresetdone_i)
    begin
        if(gt3_rxresetdone_i = '0') then
            gt3_rxresetdone_r  <= '0'   after DLY;
            gt3_rxresetdone_r2 <= '0'   after DLY;
        elsif(gt3_rxusrclk_i'event and gt3_rxusrclk_i = '1') then
            gt3_rxresetdone_r  <= gt3_rxresetdone_i   after DLY;
            gt3_rxresetdone_r2 <= gt3_rxresetdone_r   after DLY;
            gt3_rxresetdone_r3  <= gt3_rxresetdone_r2   after DLY;
        end if;
    end process;


    process( gt0_txusrclk_i,gt3_txfsmresetdone_i)
    begin
        if(gt3_txfsmresetdone_i = '0') then
            gt3_txfsmresetdone_r  <= '0'   after DLY;
            gt3_txfsmresetdone_r2 <= '0'   after DLY;
        elsif(gt0_txusrclk_i'event and gt0_txusrclk_i = '1') then
            gt3_txfsmresetdone_r  <= gt3_txfsmresetdone_i   after DLY;
            gt3_txfsmresetdone_r2 <= gt3_txfsmresetdone_r   after DLY;
        end if;
    end process;

    ------------------------------ Frame Generators ---------------------------
    -- The example design uses Block RAM based frame generators to provide test
    -- data to the GTs for transmission. By default the frame generators are 
    -- loaded with an incrementing data sequence that includes commas/alignment
    -- characters for alignment. If your protocol uses channel bonding, the 
    -- frame generator will also be preloaded with a channel bonding sequence.
    
    -- You can modify the data transmitted by changing the INIT values of the frame
    -- generator in this file. Pay careful attention to bit order and the spacing
    -- of your control and alignment characters.

    gt0_frame_gen : xilinx_gth_16b_5g_cpll_GT_FRAME_GEN
    generic map
    (
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM
    )
    port map
    (
        -- User Interface
        TX_DATA_OUT(79 downto 32)       =>      gt0_txdata_float_i,
        TX_DATA_OUT(15 downto 0)        =>      gt0_txdata_float16_i,
        TX_DATA_OUT(31 downto 16)       =>      gt0_txdata_i,
 
        TXCTRL_OUT(7 downto 2)          =>      gt0_txcharisk_float_i,
        TXCTRL_OUT(1 downto 0)          =>      gt0_txcharisk_i,
        -- System Interface
        USER_CLK                        =>      gt0_txusrclk_i,
        SYSTEM_RESET                    =>      gt0_tx_system_reset_c
    );
    
    gt1_frame_gen : xilinx_gth_16b_5g_cpll_GT_FRAME_GEN
    generic map
    (
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM
    )
    port map
    (
        -- User Interface
        TX_DATA_OUT(79 downto 32)       =>      gt1_txdata_float_i,
        TX_DATA_OUT(15 downto 0)        =>      gt1_txdata_float16_i,
        TX_DATA_OUT(31 downto 16)       =>      gt1_txdata_i,
 
        TXCTRL_OUT(7 downto 2)          =>      gt1_txcharisk_float_i,
        TXCTRL_OUT(1 downto 0)          =>      gt1_txcharisk_i,
        -- System Interface
        USER_CLK                        =>      gt0_txusrclk_i,
        SYSTEM_RESET                    =>      gt1_tx_system_reset_c
    );
    
    gt2_frame_gen : xilinx_gth_16b_5g_cpll_GT_FRAME_GEN
    generic map
    (
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM
    )
    port map
    (
        -- User Interface
        TX_DATA_OUT(79 downto 32)       =>      gt2_txdata_float_i,
        TX_DATA_OUT(15 downto 0)        =>      gt2_txdata_float16_i,
        TX_DATA_OUT(31 downto 16)       =>      gt2_txdata_i,
 
        TXCTRL_OUT(7 downto 2)          =>      gt2_txcharisk_float_i,
        TXCTRL_OUT(1 downto 0)          =>      gt2_txcharisk_i,
        -- System Interface
        USER_CLK                        =>      gt0_txusrclk_i,
        SYSTEM_RESET                    =>      gt2_tx_system_reset_c
    );
    
    gt3_frame_gen : xilinx_gth_16b_5g_cpll_GT_FRAME_GEN
    generic map
    (
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM
    )
    port map
    (
        -- User Interface
        TX_DATA_OUT(79 downto 32)       =>      gt3_txdata_float_i,
        TX_DATA_OUT(15 downto 0)        =>      gt3_txdata_float16_i,
        TX_DATA_OUT(31 downto 16)       =>      gt3_txdata_i,
 
        TXCTRL_OUT(7 downto 2)          =>      gt3_txcharisk_float_i,
        TXCTRL_OUT(1 downto 0)          =>      gt3_txcharisk_i,
        -- System Interface
        USER_CLK                        =>      gt0_txusrclk_i,
        SYSTEM_RESET                    =>      gt3_tx_system_reset_c
    );
    


    ---------------------------------- Frame Checkers -------------------------
    -- The example design uses Block RAM based frame checkers to verify incoming  
    -- data. By default the frame generators are loaded with a data sequence that 
    -- matches the outgoing sequence of the frame generators for the TX ports.
    
    -- You can modify the expected data sequence by changing the INIT values of the frame
    -- checkers in this file. Pay careful attention to bit order and the spacing
    -- of your control and alignment characters.
    
    -- When the frame checker receives data, it attempts to synchronise to the 
    -- incoming pattern by looking for the first sequence in the pattern. Once it 
    -- finds the first sequence, it increments through the sequence, and indicates an 
    -- error whenever the next value received does not match the expected value.

    gt0_frame_check_reset_i                      <= reset_on_data_error_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else gt0_matchn_i;

    -- gt0_frame_check0 is always connected to the lane with the start of char
    -- and this lane starts off the data checking on all the other lanes. The INC_IN port is tied off
    gt0_inc_in_i                                 <= '0';

    gt0_frame_check : xilinx_gth_16b_5g_cpll_GT_FRAME_CHECK
    generic map
    (
        RX_DATA_WIDTH                   =>      16,
        RXCTRL_WIDTH                    =>      2,
        COMMA_DOUBLE                    =>      x"02bc",
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        START_OF_PACKET_CHAR            =>      x"02bc"
    )
    port map
    (
        -- GT Interface
        RX_DATA_IN                      =>      gt0_rxdata_i,
        RXCTRL_IN                       =>      gt0_rxcharisk_i,
        RXENMCOMMADET_OUT               =>      gt0_rxmcommaalignen_i,
        RXENPCOMMADET_OUT               =>      gt0_rxpcommaalignen_i,
        RX_ENCHAN_SYNC_OUT              =>      open,
        RX_CHANBOND_SEQ_IN              =>      tied_to_ground_i,
        -- Control Interface
        INC_IN                          =>      gt0_inc_in_i,
        INC_OUT                         =>      gt0_inc_out_i,
        PATTERN_MATCHB_OUT              =>      gt0_matchn_i,
        RESET_ON_ERROR_IN               =>      gt0_frame_check_reset_i,
        -- System Interface
        USER_CLK                        =>      gt0_rxusrclk_i,
        SYSTEM_RESET                    =>      gt0_rx_system_reset_c,
        ERROR_COUNT_OUT                 =>      gt0_error_count_i,
        TRACK_DATA_OUT                  =>      gt0_track_data_i
    );

    gt1_frame_check_reset_i                      <= reset_on_data_error_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else gt1_matchn_i;

    -- in the "independent lanes" configuration, each of the lanes looks for the unique start char and
    -- in this case, the INC_IN port is tied off.
    -- Else, the data checking is triggered by the "master" lane
    gt1_inc_in_i                                 <= gt0_inc_out_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else '0';

    gt1_frame_check : xilinx_gth_16b_5g_cpll_GT_FRAME_CHECK
    generic map
    (
        RX_DATA_WIDTH                   =>      16,
        RXCTRL_WIDTH                    =>      2,
        COMMA_DOUBLE                    =>      x"02bc",
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        START_OF_PACKET_CHAR            =>      x"02bc"
    )
    port map
    (
        -- GT Interface
        RX_DATA_IN                      =>      gt1_rxdata_i,
        RXCTRL_IN                       =>      gt1_rxcharisk_i,
        RXENMCOMMADET_OUT               =>      gt1_rxmcommaalignen_i,
        RXENPCOMMADET_OUT               =>      gt1_rxpcommaalignen_i,
        RX_ENCHAN_SYNC_OUT              =>      open,
        RX_CHANBOND_SEQ_IN              =>      tied_to_ground_i,
        -- Control Interface
        INC_IN                          =>      gt1_inc_in_i,
        INC_OUT                         =>      gt1_inc_out_i,
        PATTERN_MATCHB_OUT              =>      gt1_matchn_i,
        RESET_ON_ERROR_IN               =>      gt1_frame_check_reset_i,
        -- System Interface
        USER_CLK                        =>      gt1_rxusrclk_i,
        SYSTEM_RESET                    =>      gt1_rx_system_reset_c,
        ERROR_COUNT_OUT                 =>      gt1_error_count_i,
        TRACK_DATA_OUT                  =>      gt1_track_data_i
    );

    gt2_frame_check_reset_i                      <= reset_on_data_error_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else gt2_matchn_i;

    -- in the "independent lanes" configuration, each of the lanes looks for the unique start char and
    -- in this case, the INC_IN port is tied off.
    -- Else, the data checking is triggered by the "master" lane
    gt2_inc_in_i                                 <= gt0_inc_out_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else '0';

    gt2_frame_check : xilinx_gth_16b_5g_cpll_GT_FRAME_CHECK
    generic map
    (
        RX_DATA_WIDTH                   =>      16,
        RXCTRL_WIDTH                    =>      2,
        COMMA_DOUBLE                    =>      x"02bc",
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        START_OF_PACKET_CHAR            =>      x"02bc"
    )
    port map
    (
        -- GT Interface
        RX_DATA_IN                      =>      gt2_rxdata_i,
        RXCTRL_IN                       =>      gt2_rxcharisk_i,
        RXENMCOMMADET_OUT               =>      gt2_rxmcommaalignen_i,
        RXENPCOMMADET_OUT               =>      gt2_rxpcommaalignen_i,
        RX_ENCHAN_SYNC_OUT              =>      open,
        RX_CHANBOND_SEQ_IN              =>      tied_to_ground_i,
        -- Control Interface
        INC_IN                          =>      gt2_inc_in_i,
        INC_OUT                         =>      gt2_inc_out_i,
        PATTERN_MATCHB_OUT              =>      gt2_matchn_i,
        RESET_ON_ERROR_IN               =>      gt2_frame_check_reset_i,
        -- System Interface
        USER_CLK                        =>      gt2_rxusrclk_i,
        SYSTEM_RESET                    =>      gt2_rx_system_reset_c,
        ERROR_COUNT_OUT                 =>      gt2_error_count_i,
        TRACK_DATA_OUT                  =>      gt2_track_data_i
    );

    gt3_frame_check_reset_i                      <= reset_on_data_error_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else gt3_matchn_i;

    -- in the "independent lanes" configuration, each of the lanes looks for the unique start char and
    -- in this case, the INC_IN port is tied off.
    -- Else, the data checking is triggered by the "master" lane
    gt3_inc_in_i                                 <= gt0_inc_out_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else '0';

    gt3_frame_check : xilinx_gth_16b_5g_cpll_GT_FRAME_CHECK
    generic map
    (
        RX_DATA_WIDTH                   =>      16,
        RXCTRL_WIDTH                    =>      2,
        COMMA_DOUBLE                    =>      x"02bc",
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        START_OF_PACKET_CHAR            =>      x"02bc"
    )
    port map
    (
        -- GT Interface
        RX_DATA_IN                      =>      gt3_rxdata_i,
        RXCTRL_IN                       =>      gt3_rxcharisk_i,
        RXENMCOMMADET_OUT               =>      gt3_rxmcommaalignen_i,
        RXENPCOMMADET_OUT               =>      gt3_rxpcommaalignen_i,
        RX_ENCHAN_SYNC_OUT              =>      open,
        RX_CHANBOND_SEQ_IN              =>      tied_to_ground_i,
        -- Control Interface
        INC_IN                          =>      gt3_inc_in_i,
        INC_OUT                         =>      gt3_inc_out_i,
        PATTERN_MATCHB_OUT              =>      gt3_matchn_i,
        RESET_ON_ERROR_IN               =>      gt3_frame_check_reset_i,
        -- System Interface
        USER_CLK                        =>      gt3_rxusrclk_i,
        SYSTEM_RESET                    =>      gt3_rx_system_reset_c,
        ERROR_COUNT_OUT                 =>      gt3_error_count_i,
        TRACK_DATA_OUT                  =>      gt3_track_data_i
    );




    TRACK_DATA_OUT                               <= track_data_out_i;

    track_data_out_i                             <= 
                                gt0_track_data_i  and
                                gt1_track_data_i  and
                                gt2_track_data_i  and
                                gt3_track_data_i ;














-------------------------------------------------------------------------------
    
    
    
    
    

----------------------------- Chipscope Connections -----------------------
    -- When the example design is run in hardware, it uses chipscope to allow the
    -- example design and GT wrapper to be controlled and monitored. The 
    -- EXAMPLE_USE_CHIPSCOPE parameter allows chipscope to be removed for simulation.

chipscope : if EXAMPLE_USE_CHIPSCOPE = 1 generate
    
    -- ICON for all VIOs 
    icon_i : icon
    port map
    (
        control0                        =>      shared_vio_control_i,
        control1                        =>      tx_data_vio_control_i,
        control2                        =>      rx_data_vio_control_i,
        control3                        =>      ila_control_i,
        control4                        =>      channel_drp_vio_control_i,
        control5                        =>      common_drp_vio_control_i
    );

    -- Shared VIO for Channel DRP  
    channel_drp_i : data_vio 
    port map
    (
        control                         =>      channel_drp_vio_control_i,
        async_in                        =>      channel_drp_vio_async_in_i,
        async_out                       =>      channel_drp_vio_async_out_i,
        sync_in                         =>      channel_drp_vio_sync_in_i,
        sync_out                        =>      channel_drp_vio_sync_out_i,
        clk                             =>      drpclk_in_i
    );

    -- Shared VIO for Quad common DRP  
    common_drp_i : data_vio 
    port map
    (
        control                         =>      common_drp_vio_control_i,
        async_in                        =>      common_drp_vio_async_in_i,
        async_out                       =>      common_drp_vio_async_out_i,
        sync_in                         =>      common_drp_vio_sync_in_i,
        sync_out                        =>      common_drp_vio_sync_out_i,
        clk                             =>      drpclk_in_i
    );

    -- Shared VIO for all transievers 
    shared_vio_i : data_vio
    port map
    (
        control                         =>      shared_vio_control_i,
        clk                             =>      tied_to_ground_i,
        async_in                        =>      shared_vio_in_i,
        async_out                       =>      shared_vio_out_i,
        sync_in                         =>      tied_to_ground_vec_i(31 downto 0),
        sync_out                        =>      open
    );
    
    
    -- TX VIO 
    tx_data_vio_i : data_vio
    port map
    (
        control                         =>      tx_data_vio_control_i,
        clk                             =>      gt0_txusrclk_i,
        async_in                        =>      tx_data_vio_async_in_i,
        async_out                       =>      tx_data_vio_async_out_i,
        sync_in                         =>      tx_data_vio_sync_in_i,
        sync_out                        =>      tx_data_vio_sync_out_i
    );
    
    -- RX VIO 
    rx_data_vio_i : data_vio
    port map
    (
        control                         =>      rx_data_vio_control_i,
        clk                             =>      rx_vio_ila_clk_i,
        async_in                        =>      rx_data_vio_async_in_i,
        async_out                       =>      rx_data_vio_async_out_i,
        sync_in                         =>      rx_data_vio_sync_in_i,
        sync_out                        =>      rx_data_vio_sync_out_i
    );
    
    -- RX ILA
    ila_i : ila
    port map
    (
        control                         =>      ila_control_i,
        clk                             =>      rx_vio_ila_clk_i,
        trig0                           =>      ila_in_i
    );


    -- The RX VIO and ILA uses GT0's RXUSRCLK2
    rx_vio_ila_clk_i <= gt0_rxusrclk_i;

    -- assign resets for frame_gen modules

    gt0_tx_system_reset_c                        <= not gt0_txfsmresetdone_r2 or user_tx_reset_i;

    gt1_tx_system_reset_c                        <= not gt1_txfsmresetdone_r2 or user_tx_reset_i;

    gt2_tx_system_reset_c                        <= not gt2_txfsmresetdone_r2 or user_tx_reset_i;

    gt3_tx_system_reset_c                        <= not gt3_txfsmresetdone_r2 or user_tx_reset_i;

    -- assign resets for frame_check modules
    gt0_rx_system_reset_c                        <= not gt0_rxresetdone_r3 or user_rx_reset_i;
    gt1_rx_system_reset_c                        <= not gt1_rxresetdone_r3 or user_rx_reset_i;
    gt2_rx_system_reset_c                        <= not gt2_rxresetdone_r3 or user_rx_reset_i;
    gt3_rx_system_reset_c                        <= not gt3_rxresetdone_r3 or user_rx_reset_i;

    gt0_gtrxreset_i                              <= gtrxreset_i or not gt0_cplllock_i;
    gt0_gttxreset_i                              <= gttxreset_i or not gt0_cplllock_i;
    gt1_gtrxreset_i                              <= gtrxreset_i or not gt1_cplllock_i;
    gt1_gttxreset_i                              <= gttxreset_i or not gt1_cplllock_i;
    gt2_gtrxreset_i                              <= gtrxreset_i or not gt2_cplllock_i;
    gt2_gttxreset_i                              <= gttxreset_i or not gt2_cplllock_i;
    gt3_gtrxreset_i                              <= gtrxreset_i or not gt3_cplllock_i;
    gt3_gttxreset_i                              <= gttxreset_i or not gt3_cplllock_i;

    gt0_cpllreset_i                              <= cpllreset_i;
    gt1_cpllreset_i                              <= cpllreset_i;
    gt2_cpllreset_i                              <= cpllreset_i;
    gt3_cpllreset_i                              <= cpllreset_i;


    -- Shared VIO Outputs
    gttxreset_i                                  <= shared_vio_out_i(31);
    gtrxreset_i                                  <= shared_vio_out_i(30);
    user_tx_reset_i                              <= shared_vio_out_i(29);
    user_rx_reset_i                              <= shared_vio_out_i(28);
    mux_sel_i                                    <= shared_vio_out_i(27 downto 26);
    cpllreset_i                                  <= shared_vio_out_i(25);

    -- Shared VIO Inputs
    shared_vio_in_i(31 downto 0)                 <= "00000000000000000000000000000000";

    -- Chipscope connections on GT 0
    gt0_tx_data_vio_async_in_i(31 downto 0)      <= "00000000000000000000000000000000";
    gt0_tx_data_vio_sync_in_i(31)                <= gt0_txresetdone_i;
    gt0_tx_data_vio_sync_in_i(30 downto 0)       <= "0000000000000000000000000000000";
    gt0_loopback_i                               <= tx_data_vio_async_out_i(31 downto 29);
    gt0_txuserrdy_i                              <= tx_data_vio_sync_out_i(31);
    gt0_txprbssel_i                              <= tx_data_vio_sync_out_i(30 downto 28);
    gt0_txpolarity_i                             <= tx_data_vio_sync_out_i(27);
    gt0_rx_data_vio_async_in_i(31 downto 0)      <= "00000000000000000000000000000000";
    gt0_rx_data_vio_sync_in_i(31)                <= gt0_rxresetdone_i;
    gt0_rx_data_vio_sync_in_i(30 downto 0)       <= "0000000000000000000000000000000";
    gt0_rxuserrdy_i                              <= rx_data_vio_async_out_i(31);
    gt0_rxprbscntreset_i                         <= rx_data_vio_sync_out_i(31);
    gt0_rxprbssel_i                              <= rx_data_vio_sync_out_i(30 downto 28);
    gt0_rxpolarity_i                             <= rx_data_vio_sync_out_i(27);
    gt0_ila_in_i(163 downto 162)                 <= gt0_rxchariscomma_i;
    gt0_ila_in_i(161 downto 160)                 <= gt0_rxcharisk_i;
    gt0_ila_in_i(159 downto 158)                 <= gt0_rxdisperr_i;
    gt0_ila_in_i(157 downto 156)                 <= gt0_rxnotintable_i;
    gt0_ila_in_i(155)                            <= gt0_rxbyteisaligned_i;
    gt0_ila_in_i(154)                            <= gt0_rxcommadet_i;
    gt0_ila_in_i(153)                            <= gt0_rxprbserr_i;
    gt0_ila_in_i(152 downto 137)                 <= gt0_rxdata_i;
    gt0_ila_in_i(136 downto 129)                 <= gt0_error_count_i;
    gt0_ila_in_i(128)                            <= gt0_track_data_i;
    gt0_ila_in_i(127 downto 0)                   <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    gt0_channel_drp_vio_async_in_i(31)           <= gt0_drprdy_i;
    gt0_channel_drp_vio_async_in_i(30 downto 15) <= gt0_drpdo_i;
    gt0_channel_drp_vio_async_in_i(14 downto 0)  <= "000000000000000";
    gt0_channel_drp_vio_sync_in_i(31 downto 0)   <= "00000000000000000000000000000000";
    gt0_drpaddr_i                                <= channel_drp_vio_async_out_i(31 downto 23);
    gt0_drpdi_i                                  <= channel_drp_vio_async_out_i(22 downto 7);
    gt0_drpen_i                                  <= channel_drp_vio_async_out_i(6);
    gt0_drpwe_i                                  <= channel_drp_vio_async_out_i(5);
    gt0_common_drp_vio_async_in_i(31 downto 0)   <= "00000000000000000000000000000000";
    gt0_common_drp_vio_sync_in_i(31 downto 0)    <= "00000000000000000000000000000000";

    -- Chipscope connections on GT 1
    gt1_tx_data_vio_async_in_i(31 downto 0)      <= "00000000000000000000000000000000";
    gt1_tx_data_vio_sync_in_i(31)                <= gt1_txresetdone_i;
    gt1_tx_data_vio_sync_in_i(30 downto 0)       <= "0000000000000000000000000000000";
    gt1_loopback_i                               <= tx_data_vio_async_out_i(31 downto 29);
    gt1_txuserrdy_i                              <= tx_data_vio_sync_out_i(31);
    gt1_txprbssel_i                              <= tx_data_vio_sync_out_i(30 downto 28);
    gt1_txpolarity_i                             <= tx_data_vio_sync_out_i(27);
    gt1_rx_data_vio_async_in_i(31 downto 0)      <= "00000000000000000000000000000000";
    gt1_rx_data_vio_sync_in_i(31)                <= gt1_rxresetdone_i;
    gt1_rx_data_vio_sync_in_i(30 downto 0)       <= "0000000000000000000000000000000";
    gt1_rxuserrdy_i                              <= rx_data_vio_async_out_i(31);
    gt1_rxprbscntreset_i                         <= rx_data_vio_sync_out_i(31);
    gt1_rxprbssel_i                              <= rx_data_vio_sync_out_i(30 downto 28);
    gt1_rxpolarity_i                             <= rx_data_vio_sync_out_i(27);
    gt1_ila_in_i(163 downto 162)                 <= gt1_rxchariscomma_i;
    gt1_ila_in_i(161 downto 160)                 <= gt1_rxcharisk_i;
    gt1_ila_in_i(159 downto 158)                 <= gt1_rxdisperr_i;
    gt1_ila_in_i(157 downto 156)                 <= gt1_rxnotintable_i;
    gt1_ila_in_i(155)                            <= gt1_rxbyteisaligned_i;
    gt1_ila_in_i(154)                            <= gt1_rxcommadet_i;
    gt1_ila_in_i(153)                            <= gt1_rxprbserr_i;
    gt1_ila_in_i(152 downto 137)                 <= gt1_rxdata_i;
    gt1_ila_in_i(136 downto 129)                 <= gt1_error_count_i;
    gt1_ila_in_i(128)                            <= gt1_track_data_i;
    gt1_ila_in_i(127 downto 0)                   <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    gt1_channel_drp_vio_async_in_i(31)           <= gt1_drprdy_i;
    gt1_channel_drp_vio_async_in_i(30 downto 15) <= gt1_drpdo_i;
    gt1_channel_drp_vio_async_in_i(14 downto 0)  <= "000000000000000";
    gt1_channel_drp_vio_sync_in_i(31 downto 0)   <= "00000000000000000000000000000000";
    gt1_drpaddr_i                                <= channel_drp_vio_async_out_i(31 downto 23);
    gt1_drpdi_i                                  <= channel_drp_vio_async_out_i(22 downto 7);
    gt1_drpen_i                                  <= channel_drp_vio_async_out_i(6);
    gt1_drpwe_i                                  <= channel_drp_vio_async_out_i(5);

    -- Chipscope connections on GT 2
    gt2_tx_data_vio_async_in_i(31 downto 0)      <= "00000000000000000000000000000000";
    gt2_tx_data_vio_sync_in_i(31)                <= gt2_txresetdone_i;
    gt2_tx_data_vio_sync_in_i(30 downto 0)       <= "0000000000000000000000000000000";
    gt2_loopback_i                               <= tx_data_vio_async_out_i(31 downto 29);
    gt2_txuserrdy_i                              <= tx_data_vio_sync_out_i(31);
    gt2_txprbssel_i                              <= tx_data_vio_sync_out_i(30 downto 28);
    gt2_txpolarity_i                             <= tx_data_vio_sync_out_i(27);
    gt2_rx_data_vio_async_in_i(31 downto 0)      <= "00000000000000000000000000000000";
    gt2_rx_data_vio_sync_in_i(31)                <= gt2_rxresetdone_i;
    gt2_rx_data_vio_sync_in_i(30 downto 0)       <= "0000000000000000000000000000000";
    gt2_rxuserrdy_i                              <= rx_data_vio_async_out_i(31);
    gt2_rxprbscntreset_i                         <= rx_data_vio_sync_out_i(31);
    gt2_rxprbssel_i                              <= rx_data_vio_sync_out_i(30 downto 28);
    gt2_rxpolarity_i                             <= rx_data_vio_sync_out_i(27);
    gt2_ila_in_i(163 downto 162)                 <= gt2_rxchariscomma_i;
    gt2_ila_in_i(161 downto 160)                 <= gt2_rxcharisk_i;
    gt2_ila_in_i(159 downto 158)                 <= gt2_rxdisperr_i;
    gt2_ila_in_i(157 downto 156)                 <= gt2_rxnotintable_i;
    gt2_ila_in_i(155)                            <= gt2_rxbyteisaligned_i;
    gt2_ila_in_i(154)                            <= gt2_rxcommadet_i;
    gt2_ila_in_i(153)                            <= gt2_rxprbserr_i;
    gt2_ila_in_i(152 downto 137)                 <= gt2_rxdata_i;
    gt2_ila_in_i(136 downto 129)                 <= gt2_error_count_i;
    gt2_ila_in_i(128)                            <= gt2_track_data_i;
    gt2_ila_in_i(127 downto 0)                   <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    gt2_channel_drp_vio_async_in_i(31)           <= gt2_drprdy_i;
    gt2_channel_drp_vio_async_in_i(30 downto 15) <= gt2_drpdo_i;
    gt2_channel_drp_vio_async_in_i(14 downto 0)  <= "000000000000000";
    gt2_channel_drp_vio_sync_in_i(31 downto 0)   <= "00000000000000000000000000000000";
    gt2_drpaddr_i                                <= channel_drp_vio_async_out_i(31 downto 23);
    gt2_drpdi_i                                  <= channel_drp_vio_async_out_i(22 downto 7);
    gt2_drpen_i                                  <= channel_drp_vio_async_out_i(6);
    gt2_drpwe_i                                  <= channel_drp_vio_async_out_i(5);

    -- Chipscope connections on GT 3
    gt3_tx_data_vio_async_in_i(31 downto 0)      <= "00000000000000000000000000000000";
    gt3_tx_data_vio_sync_in_i(31)                <= gt3_txresetdone_i;
    gt3_tx_data_vio_sync_in_i(30 downto 0)       <= "0000000000000000000000000000000";
    gt3_loopback_i                               <= tx_data_vio_async_out_i(31 downto 29);
    gt3_txuserrdy_i                              <= tx_data_vio_sync_out_i(31);
    gt3_txprbssel_i                              <= tx_data_vio_sync_out_i(30 downto 28);
    gt3_txpolarity_i                             <= tx_data_vio_sync_out_i(27);
    gt3_rx_data_vio_async_in_i(31 downto 0)      <= "00000000000000000000000000000000";
    gt3_rx_data_vio_sync_in_i(31)                <= gt3_rxresetdone_i;
    gt3_rx_data_vio_sync_in_i(30 downto 0)       <= "0000000000000000000000000000000";
    gt3_rxuserrdy_i                              <= rx_data_vio_async_out_i(31);
    gt3_rxprbscntreset_i                         <= rx_data_vio_sync_out_i(31);
    gt3_rxprbssel_i                              <= rx_data_vio_sync_out_i(30 downto 28);
    gt3_rxpolarity_i                             <= rx_data_vio_sync_out_i(27);
    gt3_ila_in_i(163 downto 162)                 <= gt3_rxchariscomma_i;
    gt3_ila_in_i(161 downto 160)                 <= gt3_rxcharisk_i;
    gt3_ila_in_i(159 downto 158)                 <= gt3_rxdisperr_i;
    gt3_ila_in_i(157 downto 156)                 <= gt3_rxnotintable_i;
    gt3_ila_in_i(155)                            <= gt3_rxbyteisaligned_i;
    gt3_ila_in_i(154)                            <= gt3_rxcommadet_i;
    gt3_ila_in_i(153)                            <= gt3_rxprbserr_i;
    gt3_ila_in_i(152 downto 137)                 <= gt3_rxdata_i;
    gt3_ila_in_i(136 downto 129)                 <= gt3_error_count_i;
    gt3_ila_in_i(128)                            <= gt3_track_data_i;
    gt3_ila_in_i(127 downto 0)                   <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    gt3_channel_drp_vio_async_in_i(31)           <= gt3_drprdy_i;
    gt3_channel_drp_vio_async_in_i(30 downto 15) <= gt3_drpdo_i;
    gt3_channel_drp_vio_async_in_i(14 downto 0)  <= "000000000000000";
    gt3_channel_drp_vio_sync_in_i(31 downto 0)   <= "00000000000000000000000000000000";
    gt3_drpaddr_i                                <= channel_drp_vio_async_out_i(31 downto 23);
    gt3_drpdi_i                                  <= channel_drp_vio_async_out_i(22 downto 7);
    gt3_drpen_i                                  <= channel_drp_vio_async_out_i(6);
    gt3_drpwe_i                                  <= channel_drp_vio_async_out_i(5);


    tx_data_vio_async_in_i              <=      gt0_tx_data_vio_async_in_i when (mux_sel_i = "00")
                                        else    gt1_tx_data_vio_async_in_i when (mux_sel_i = "01")
                                        else    gt2_tx_data_vio_async_in_i when (mux_sel_i = "10")
                                        else    gt3_tx_data_vio_async_in_i;

    tx_data_vio_sync_in_i               <=      gt0_tx_data_vio_sync_in_i when (mux_sel_i = "00")
                                        else    gt1_tx_data_vio_sync_in_i when (mux_sel_i = "01")
                                        else    gt2_tx_data_vio_sync_in_i when (mux_sel_i = "10")
                                        else    gt3_tx_data_vio_sync_in_i;


    rx_data_vio_async_in_i              <=      gt0_rx_data_vio_async_in_i when (mux_sel_i = "00")
                                        else    gt1_rx_data_vio_async_in_i when (mux_sel_i = "01")
                                        else    gt2_rx_data_vio_async_in_i when (mux_sel_i = "10")
                                        else    gt3_rx_data_vio_async_in_i;

    rx_data_vio_sync_in_i               <=      gt0_rx_data_vio_sync_in_i when (mux_sel_i = "00")
                                        else    gt1_rx_data_vio_sync_in_i when (mux_sel_i = "01")
                                        else    gt2_rx_data_vio_sync_in_i when (mux_sel_i = "10")
                                        else    gt3_rx_data_vio_sync_in_i;

    ila_in_i                            <=      gt0_ila_in_i when (mux_sel_i = "00")
                                        else    gt1_ila_in_i when (mux_sel_i = "01")
                                        else    gt2_ila_in_i when (mux_sel_i = "10")
                                        else    gt3_ila_in_i;


    channel_drp_vio_async_in_i          <=      gt0_channel_drp_vio_async_in_i when (mux_sel_i = "00")
                                        else    gt1_channel_drp_vio_async_in_i when (mux_sel_i = "01")
                                        else    gt2_channel_drp_vio_async_in_i when (mux_sel_i = "10")
                                        else    gt3_channel_drp_vio_async_in_i;

    channel_drp_vio_sync_in_i           <=      gt0_channel_drp_vio_sync_in_i when (mux_sel_i = "00")
                                        else    gt1_channel_drp_vio_sync_in_i when (mux_sel_i = "01")
                                        else    gt2_channel_drp_vio_sync_in_i when (mux_sel_i = "10")
                                        else    gt3_channel_drp_vio_sync_in_i;

    common_drp_vio_async_in_i <= (others => '0');
    common_drp_vio_sync_in_i  <= (others => '0');

end generate chipscope;

no_chipscope : if EXAMPLE_USE_CHIPSCOPE = 0 generate


    -- assign resets for frame_gen modules
    gt0_tx_system_reset_c                        <= not gt0_txfsmresetdone_r2;
    gt1_tx_system_reset_c                        <= not gt1_txfsmresetdone_r2;
    gt2_tx_system_reset_c                        <= not gt2_txfsmresetdone_r2;
    gt3_tx_system_reset_c                        <= not gt3_txfsmresetdone_r2;

    -- assign resets for frame_check modules
    gt0_rx_system_reset_c                        <= not gt0_rxresetdone_r3;
    gt1_rx_system_reset_c                        <= not gt1_rxresetdone_r3;
    gt2_rx_system_reset_c                        <= not gt2_rxresetdone_r3;
    gt3_rx_system_reset_c                        <= not gt3_rxresetdone_r3;

    gttxreset_i                                  <= tied_to_ground_i;
    gtrxreset_i                                  <= tied_to_ground_i;
    user_tx_reset_i                              <= tied_to_ground_i;
    user_rx_reset_i                              <= tied_to_ground_i;
    mux_sel_i                                    <= tied_to_ground_vec_i(1 downto 0);
    gt0_loopback_i                               <= tied_to_ground_vec_i(2 downto 0);
    gt0_txprbssel_i                              <= tied_to_ground_vec_i(2 downto 0);
    gt0_txpolarity_i                             <= tied_to_ground_i;
    gt0_rxprbscntreset_i                         <= tied_to_ground_i;
    gt0_rxprbssel_i                              <= tied_to_ground_vec_i(2 downto 0);
    gt0_rxpolarity_i                             <= tied_to_ground_i;
    gt0_drpaddr_i                                <= tied_to_ground_vec_i(8 downto 0);
    gt0_drpdi_i                                  <= tied_to_ground_vec_i(15 downto 0);
    gt0_drpen_i                                  <= tied_to_ground_i;
    gt0_drpwe_i                                  <= tied_to_ground_i;
    gt1_loopback_i                               <= tied_to_ground_vec_i(2 downto 0);
    gt1_txprbssel_i                              <= tied_to_ground_vec_i(2 downto 0);
    gt1_txpolarity_i                             <= tied_to_ground_i;
    gt1_rxprbscntreset_i                         <= tied_to_ground_i;
    gt1_rxprbssel_i                              <= tied_to_ground_vec_i(2 downto 0);
    gt1_rxpolarity_i                             <= tied_to_ground_i;
    gt1_drpaddr_i                                <= tied_to_ground_vec_i(8 downto 0);
    gt1_drpdi_i                                  <= tied_to_ground_vec_i(15 downto 0);
    gt1_drpen_i                                  <= tied_to_ground_i;
    gt1_drpwe_i                                  <= tied_to_ground_i;
    gt2_loopback_i                               <= tied_to_ground_vec_i(2 downto 0);
    gt2_txprbssel_i                              <= tied_to_ground_vec_i(2 downto 0);
    gt2_txpolarity_i                             <= tied_to_ground_i;
    gt2_rxprbscntreset_i                         <= tied_to_ground_i;
    gt2_rxprbssel_i                              <= tied_to_ground_vec_i(2 downto 0);
    gt2_rxpolarity_i                             <= tied_to_ground_i;
    gt2_drpaddr_i                                <= tied_to_ground_vec_i(8 downto 0);
    gt2_drpdi_i                                  <= tied_to_ground_vec_i(15 downto 0);
    gt2_drpen_i                                  <= tied_to_ground_i;
    gt2_drpwe_i                                  <= tied_to_ground_i;
    gt3_loopback_i                               <= tied_to_ground_vec_i(2 downto 0);
    gt3_txprbssel_i                              <= tied_to_ground_vec_i(2 downto 0);
    gt3_txpolarity_i                             <= tied_to_ground_i;
    gt3_rxprbscntreset_i                         <= tied_to_ground_i;
    gt3_rxprbssel_i                              <= tied_to_ground_vec_i(2 downto 0);
    gt3_rxpolarity_i                             <= tied_to_ground_i;
    gt3_drpaddr_i                                <= tied_to_ground_vec_i(8 downto 0);
    gt3_drpdi_i                                  <= tied_to_ground_vec_i(15 downto 0);
    gt3_drpen_i                                  <= tied_to_ground_i;
    gt3_drpwe_i                                  <= tied_to_ground_i;


end generate no_chipscope;
end RTL;


