
library IEEE;
use IEEE.STD_LOGIC_1164.all;


package hgc_constants is

  constant nWafersInPanel : natural := 6;
  constant numberOfTriggerCellsPerEdge_high : natural := 5;
  constant numberOfTriggerCellsPerEdge_low  : natural := 4;
  
end hgc_constants;
